//
//    Copyright (c) 2015 Jan Adelsbach <jan@janadelsbach.com>.  
//    All Rights Reserved.
//
//    This program is free software: you can redistribute it and/or modify
//    it under the terms of the GNU General Public License as published by
//    the Free Software Foundation, either version 3 of the License, or
//    (at your option) any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program.  If not, see <http://www.gnu.org/licenses/>.
//

module mc14099b(rst, dat, wd, q);
	input rst;
	input dat;
	input wd;
	output reg [7:0] q;

	always @(rst or dat) begin
		if(rst & wd) 
			q <= 8'b0;
		else if(rst & ~wd) begin
			q    = 8'b0;
			q[a] = dat;
		end
		else if(~wd)
			q[a] <= dat;
	end
endmodule
