../../nand/nand_defines.vh