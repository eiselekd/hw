aldec/sim0/nand/nand_defines.vh