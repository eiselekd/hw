------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnologa Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=14); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

library synplify;
architecture rtl of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);
   attribute syn_ramstyle : string;
   attribute syn_ramstyle of addr_r : signal is "block_ram";

   signal ram : ram_type :=
     (
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"82c0b40c",
     3 => x"3a0b0b81",
     4 => x"bfbc0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"81c0892d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b82c0",
   162 => x"a0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8d",
   171 => x"df2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8f",
   179 => x"912d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"82c0b00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81943f82",
   257 => x"b0ac3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"ff3d0d82",
   281 => x"d0c03351",
   282 => x"70a73882",
   283 => x"c0bc0870",
   284 => x"08525270",
   285 => x"802e9438",
   286 => x"841282c0",
   287 => x"bc0c702d",
   288 => x"82c0bc08",
   289 => x"70085252",
   290 => x"70ee3881",
   291 => x"0b82d0c0",
   292 => x"34833d0d",
   293 => x"0404803d",
   294 => x"0d0b0b82",
   295 => x"d0b80880",
   296 => x"2e8e380b",
   297 => x"0b0b0b80",
   298 => x"0b802e09",
   299 => x"81068538",
   300 => x"823d0d04",
   301 => x"0b0b82d0",
   302 => x"b8510b0b",
   303 => x"0bf6c13f",
   304 => x"823d0d04",
   305 => x"04fe3d0d",
   306 => x"8d398008",
   307 => x"520b0b82",
   308 => x"b8e05189",
   309 => x"ea3f8883",
   310 => x"3f8008ee",
   311 => x"3872800c",
   312 => x"843d0d04",
   313 => x"fe3d0d82",
   314 => x"d0c40853",
   315 => x"84130870",
   316 => x"882a7081",
   317 => x"06515252",
   318 => x"70802ef0",
   319 => x"387181ff",
   320 => x"06800c84",
   321 => x"3d0d04ff",
   322 => x"3d0d82d0",
   323 => x"c4085271",
   324 => x"0870882a",
   325 => x"81327081",
   326 => x"06515151",
   327 => x"70f13873",
   328 => x"720c833d",
   329 => x"0d0482c0",
   330 => x"b008802e",
   331 => x"80c43882",
   332 => x"c0b40882",
   333 => x"2e098106",
   334 => x"9f3880c0",
   335 => x"a9808c0b",
   336 => x"82d0c40c",
   337 => x"80c0a980",
   338 => x"940b82d0",
   339 => x"c80c82b8",
   340 => x"f40b82d0",
   341 => x"bc0cb939",
   342 => x"8380800b",
   343 => x"82d0c40c",
   344 => x"82a0800b",
   345 => x"82d0c80c",
   346 => x"8290800b",
   347 => x"82d0bc0c",
   348 => x"9f39f880",
   349 => x"8080a40b",
   350 => x"82d0c40c",
   351 => x"f8808082",
   352 => x"800b82d0",
   353 => x"c80cf880",
   354 => x"8084800b",
   355 => x"82d0bc0c",
   356 => x"04f33d0d",
   357 => x"7f82d0c8",
   358 => x"08565c82",
   359 => x"750c8059",
   360 => x"805a805b",
   361 => x"7a842982",
   362 => x"d0c80805",
   363 => x"70087108",
   364 => x"719f2c7e",
   365 => x"852b5855",
   366 => x"55913df8",
   367 => x"05535957",
   368 => x"a83f7c7e",
   369 => x"7a72077c",
   370 => x"72077171",
   371 => x"60810541",
   372 => x"5f5d5b59",
   373 => x"5755817b",
   374 => x"27ca3876",
   375 => x"7c0c7784",
   376 => x"1d0c7b80",
   377 => x"0c8f3d0d",
   378 => x"048c0802",
   379 => x"8c0cf53d",
   380 => x"0d8c0894",
   381 => x"05089d38",
   382 => x"8c088c05",
   383 => x"088c0890",
   384 => x"05088c08",
   385 => x"88050858",
   386 => x"56547376",
   387 => x"0c748417",
   388 => x"0c81bf39",
   389 => x"800b8c08",
   390 => x"f0050c80",
   391 => x"0b8c08f4",
   392 => x"050c8c08",
   393 => x"8c05088c",
   394 => x"08900508",
   395 => x"5654738c",
   396 => x"08f0050c",
   397 => x"748c08f4",
   398 => x"050c8c08",
   399 => x"f8058c08",
   400 => x"f0055656",
   401 => x"88705475",
   402 => x"53765254",
   403 => x"85c13fa0",
   404 => x"0b8c0894",
   405 => x"0508318c",
   406 => x"08ec050c",
   407 => x"8c08ec05",
   408 => x"0880249d",
   409 => x"38800b8c",
   410 => x"08f4050c",
   411 => x"8c08ec05",
   412 => x"08308c08",
   413 => x"fc050871",
   414 => x"2b8c08f0",
   415 => x"050c54b9",
   416 => x"398c08fc",
   417 => x"05088c08",
   418 => x"ec05082a",
   419 => x"8c08e805",
   420 => x"0c8c08fc",
   421 => x"05088c08",
   422 => x"9405082b",
   423 => x"8c08f405",
   424 => x"0c8c08f8",
   425 => x"05088c08",
   426 => x"9405082b",
   427 => x"708c08e8",
   428 => x"0508078c",
   429 => x"08f0050c",
   430 => x"548c08f0",
   431 => x"05088c08",
   432 => x"f405088c",
   433 => x"08880508",
   434 => x"58565473",
   435 => x"760c7484",
   436 => x"170c8c08",
   437 => x"88050880",
   438 => x"0c8d3d0d",
   439 => x"8c0c048c",
   440 => x"08028c0c",
   441 => x"f93d0d80",
   442 => x"0b8c08fc",
   443 => x"050c8c08",
   444 => x"88050880",
   445 => x"25ab388c",
   446 => x"08880508",
   447 => x"308c0888",
   448 => x"050c800b",
   449 => x"8c08f405",
   450 => x"0c8c08fc",
   451 => x"05088838",
   452 => x"810b8c08",
   453 => x"f4050c8c",
   454 => x"08f40508",
   455 => x"8c08fc05",
   456 => x"0c8c088c",
   457 => x"05088025",
   458 => x"ab388c08",
   459 => x"8c050830",
   460 => x"8c088c05",
   461 => x"0c800b8c",
   462 => x"08f0050c",
   463 => x"8c08fc05",
   464 => x"08883881",
   465 => x"0b8c08f0",
   466 => x"050c8c08",
   467 => x"f005088c",
   468 => x"08fc050c",
   469 => x"80538c08",
   470 => x"8c050852",
   471 => x"8c088805",
   472 => x"085181a7",
   473 => x"3f800870",
   474 => x"8c08f805",
   475 => x"0c548c08",
   476 => x"fc050880",
   477 => x"2e8c388c",
   478 => x"08f80508",
   479 => x"308c08f8",
   480 => x"050c8c08",
   481 => x"f8050870",
   482 => x"800c5489",
   483 => x"3d0d8c0c",
   484 => x"048c0802",
   485 => x"8c0cfb3d",
   486 => x"0d800b8c",
   487 => x"08fc050c",
   488 => x"8c088805",
   489 => x"08802593",
   490 => x"388c0888",
   491 => x"0508308c",
   492 => x"0888050c",
   493 => x"810b8c08",
   494 => x"fc050c8c",
   495 => x"088c0508",
   496 => x"80258c38",
   497 => x"8c088c05",
   498 => x"08308c08",
   499 => x"8c050c81",
   500 => x"538c088c",
   501 => x"0508528c",
   502 => x"08880508",
   503 => x"51ad3f80",
   504 => x"08708c08",
   505 => x"f8050c54",
   506 => x"8c08fc05",
   507 => x"08802e8c",
   508 => x"388c08f8",
   509 => x"0508308c",
   510 => x"08f8050c",
   511 => x"8c08f805",
   512 => x"0870800c",
   513 => x"54873d0d",
   514 => x"8c0c048c",
   515 => x"08028c0c",
   516 => x"fd3d0d81",
   517 => x"0b8c08fc",
   518 => x"050c800b",
   519 => x"8c08f805",
   520 => x"0c8c088c",
   521 => x"05088c08",
   522 => x"88050827",
   523 => x"ac388c08",
   524 => x"fc050880",
   525 => x"2ea33880",
   526 => x"0b8c088c",
   527 => x"05082499",
   528 => x"388c088c",
   529 => x"0508108c",
   530 => x"088c050c",
   531 => x"8c08fc05",
   532 => x"08108c08",
   533 => x"fc050cc9",
   534 => x"398c08fc",
   535 => x"0508802e",
   536 => x"80c9388c",
   537 => x"088c0508",
   538 => x"8c088805",
   539 => x"0826a138",
   540 => x"8c088805",
   541 => x"088c088c",
   542 => x"0508318c",
   543 => x"0888050c",
   544 => x"8c08f805",
   545 => x"088c08fc",
   546 => x"0508078c",
   547 => x"08f8050c",
   548 => x"8c08fc05",
   549 => x"08812a8c",
   550 => x"08fc050c",
   551 => x"8c088c05",
   552 => x"08812a8c",
   553 => x"088c050c",
   554 => x"ffaf398c",
   555 => x"08900508",
   556 => x"802e8f38",
   557 => x"8c088805",
   558 => x"08708c08",
   559 => x"f4050c51",
   560 => x"8d398c08",
   561 => x"f8050870",
   562 => x"8c08f405",
   563 => x"0c518c08",
   564 => x"f4050880",
   565 => x"0c853d0d",
   566 => x"8c0c04fe",
   567 => x"3d0d7484",
   568 => x"1108ff11",
   569 => x"84130cff",
   570 => x"11515353",
   571 => x"80722492",
   572 => x"38720870",
   573 => x"33740881",
   574 => x"05750c80",
   575 => x"0c52843d",
   576 => x"0d047251",
   577 => x"81d83f80",
   578 => x"08800c84",
   579 => x"3d0d04fc",
   580 => x"3d0d7670",
   581 => x"797b5555",
   582 => x"55558f72",
   583 => x"278c3872",
   584 => x"75078306",
   585 => x"5170802e",
   586 => x"a738ff12",
   587 => x"5271ff2e",
   588 => x"98387270",
   589 => x"81055433",
   590 => x"74708105",
   591 => x"5634ff12",
   592 => x"5271ff2e",
   593 => x"098106ea",
   594 => x"3874800c",
   595 => x"863d0d04",
   596 => x"74517270",
   597 => x"84055408",
   598 => x"71708405",
   599 => x"530c7270",
   600 => x"84055408",
   601 => x"71708405",
   602 => x"530c7270",
   603 => x"84055408",
   604 => x"71708405",
   605 => x"530c7270",
   606 => x"84055408",
   607 => x"71708405",
   608 => x"530cf012",
   609 => x"52718f26",
   610 => x"c9388372",
   611 => x"27953872",
   612 => x"70840554",
   613 => x"08717084",
   614 => x"05530cfc",
   615 => x"12527183",
   616 => x"26ed3870",
   617 => x"54ff8339",
   618 => x"fb3d0d77",
   619 => x"893d8805",
   620 => x"55795488",
   621 => x"11085351",
   622 => x"81803f87",
   623 => x"3d0d04fc",
   624 => x"3d0d873d",
   625 => x"70708405",
   626 => x"52085653",
   627 => x"745282c0",
   628 => x"c0088811",
   629 => x"085254ab",
   630 => x"8e3f863d",
   631 => x"0d04fe3d",
   632 => x"0d747052",
   633 => x"53819fc6",
   634 => x"3fff5280",
   635 => x"08943884",
   636 => x"13081284",
   637 => x"140c7208",
   638 => x"70337408",
   639 => x"8105750c",
   640 => x"51527180",
   641 => x"0c843d0d",
   642 => x"04fd3d0d",
   643 => x"76881108",
   644 => x"5454728c",
   645 => x"38728415",
   646 => x"0c72800c",
   647 => x"853d0d04",
   648 => x"73527551",
   649 => x"80e7a03f",
   650 => x"800b8815",
   651 => x"0c800b84",
   652 => x"150c8008",
   653 => x"800c853d",
   654 => x"0d04fcc4",
   655 => x"3d0d83bf",
   656 => x"3d0883c1",
   657 => x"3d0883c3",
   658 => x"3d0883c5",
   659 => x"3d08485e",
   660 => x"484b80ee",
   661 => x"fd3f8008",
   662 => x"084c800b",
   663 => x"83bb3d0c",
   664 => x"800b83bc",
   665 => x"3d0c8070",
   666 => x"71698c05",
   667 => x"2270832a",
   668 => x"81327081",
   669 => x"06515d5d",
   670 => x"4c4f4d78",
   671 => x"6d2e0981",
   672 => x"068c3866",
   673 => x"9005086d",
   674 => x"2e098106",
   675 => x"92386651",
   676 => x"b49f3fff",
   677 => x"59800881",
   678 => x"e438668c",
   679 => x"05225a79",
   680 => x"9a065978",
   681 => x"8a2e80c0",
   682 => x"387b83a6",
   683 => x"3d707183",
   684 => x"b93d0c5e",
   685 => x"475d800b",
   686 => x"83b83d0c",
   687 => x"800b83b7",
   688 => x"3d0c8049",
   689 => x"7c5e807d",
   690 => x"337081ff",
   691 => x"065b5b5b",
   692 => x"787b2e83",
   693 => x"38815b78",
   694 => x"a52e81a9",
   695 => x"387a802e",
   696 => x"81a33881",
   697 => x"1d5ddf39",
   698 => x"668e0522",
   699 => x"70902b5a",
   700 => x"5b807924",
   701 => x"ffb33879",
   702 => x"fd065978",
   703 => x"82ba3d23",
   704 => x"7a028405",
   705 => x"89e20523",
   706 => x"669c0508",
   707 => x"82be3d0c",
   708 => x"66a40508",
   709 => x"82c03d0c",
   710 => x"b63d7082",
   711 => x"b83d0c82",
   712 => x"bb3d0c88",
   713 => x"800b82b9",
   714 => x"3d0c8880",
   715 => x"0b82bc3d",
   716 => x"0c800b82",
   717 => x"bd3d0c64",
   718 => x"537b5282",
   719 => x"b63d7052",
   720 => x"59a8a43f",
   721 => x"80085a80",
   722 => x"0b800824",
   723 => x"8f387851",
   724 => x"80d9d13f",
   725 => x"8008802e",
   726 => x"8338ff5a",
   727 => x"82b93d22",
   728 => x"70862a70",
   729 => x"8106515a",
   730 => x"5b78802e",
   731 => x"8e38668c",
   732 => x"052280c0",
   733 => x"07597867",
   734 => x"8c052379",
   735 => x"5978800c",
   736 => x"83be3d0d",
   737 => x"047c7e31",
   738 => x"5b7a802e",
   739 => x"ae387d7c",
   740 => x"0c7a841d",
   741 => x"0c83b73d",
   742 => x"081b83b8",
   743 => x"3d0c881c",
   744 => x"83b73d08",
   745 => x"811183b9",
   746 => x"3d0c8111",
   747 => x"515a5c78",
   748 => x"872480c3",
   749 => x"38681b7d",
   750 => x"335b4979",
   751 => x"81ff0659",
   752 => x"78802ea6",
   753 => x"9738811d",
   754 => x"5d807071",
   755 => x"4a4543ff",
   756 => x"416283be",
   757 => x"3d347c33",
   758 => x"5a7981ff",
   759 => x"06811e5e",
   760 => x"407fe005",
   761 => x"597880d8",
   762 => x"2686ed38",
   763 => x"78101082",
   764 => x"b9980559",
   765 => x"78080483",
   766 => x"be3ddc05",
   767 => x"526651fc",
   768 => x"883f8008",
   769 => x"89983865",
   770 => x"691c7e33",
   771 => x"5c4a5cff",
   772 => x"aa396290",
   773 => x"07436284",
   774 => x"2a708106",
   775 => x"51597898",
   776 => x"bd386286",
   777 => x"2a708106",
   778 => x"51597880",
   779 => x"2e98af38",
   780 => x"64658405",
   781 => x"8212225d",
   782 => x"4659815f",
   783 => x"800b83be",
   784 => x"3d346044",
   785 => x"80612486",
   786 => x"3862feff",
   787 => x"0643657b",
   788 => x"30707d07",
   789 => x"9f2a6630",
   790 => x"7068079f",
   791 => x"2a720752",
   792 => x"5c515b5e",
   793 => x"79802e94",
   794 => x"8c387e81",
   795 => x"2e89d538",
   796 => x"817f259a",
   797 => x"d7387e82",
   798 => x"2e8a8838",
   799 => x"82bbfc5e",
   800 => x"7d5181a2",
   801 => x"853f8008",
   802 => x"5f7e427e",
   803 => x"64258338",
   804 => x"634283bd",
   805 => x"3d337081",
   806 => x"ff065a5b",
   807 => x"78802e90",
   808 => x"90386181",
   809 => x"05426281",
   810 => x"84064160",
   811 => x"80f13867",
   812 => x"62315a80",
   813 => x"7a2580e7",
   814 => x"38907a25",
   815 => x"b43882b8",
   816 => x"f87c0c90",
   817 => x"0b841d0c",
   818 => x"83b73d08",
   819 => x"900583b8",
   820 => x"3d0c881c",
   821 => x"83b73d08",
   822 => x"811183b9",
   823 => x"3d0c8111",
   824 => x"515a5c78",
   825 => x"87248588",
   826 => x"38f01a5a",
   827 => x"799024ce",
   828 => x"3882b8f8",
   829 => x"7c0c7984",
   830 => x"1d0c83b7",
   831 => x"3d081a83",
   832 => x"b83d0c88",
   833 => x"1c83b73d",
   834 => x"08811183",
   835 => x"b93d0c81",
   836 => x"11515a5c",
   837 => x"78872492",
   838 => x"c23883bd",
   839 => x"3d335b7a",
   840 => x"81ff0659",
   841 => x"78802e8f",
   842 => x"9e3883be",
   843 => x"3dfc057c",
   844 => x"0c810b84",
   845 => x"1d0c83b7",
   846 => x"3d088105",
   847 => x"83b83d0c",
   848 => x"881c83b7",
   849 => x"3d088111",
   850 => x"83b93d0c",
   851 => x"8111515a",
   852 => x"5c788724",
   853 => x"85ec3860",
   854 => x"81802e84",
   855 => x"c338637f",
   856 => x"315a807a",
   857 => x"2580f338",
   858 => x"907a25b4",
   859 => x"3882b988",
   860 => x"7c0c900b",
   861 => x"841d0c83",
   862 => x"b73d0890",
   863 => x"0583b83d",
   864 => x"0c881c83",
   865 => x"b73d0881",
   866 => x"1183b93d",
   867 => x"0c811151",
   868 => x"5a5c7887",
   869 => x"2483f138",
   870 => x"f01a5a79",
   871 => x"9024ce38",
   872 => x"82b9887c",
   873 => x"0c79841d",
   874 => x"0c83b73d",
   875 => x"081a83b8",
   876 => x"3d0c881c",
   877 => x"83b73d08",
   878 => x"811183b9",
   879 => x"3d0c8111",
   880 => x"515a5c87",
   881 => x"79259338",
   882 => x"83be3ddc",
   883 => x"05526651",
   884 => x"f8b73f80",
   885 => x"0885c738",
   886 => x"655c6288",
   887 => x"2a813270",
   888 => x"81065159",
   889 => x"78802e8e",
   890 => x"ac387d7c",
   891 => x"0c7e841d",
   892 => x"0c83b73d",
   893 => x"081f83b8",
   894 => x"3d0c881c",
   895 => x"83b73d08",
   896 => x"811183b9",
   897 => x"3d0c8111",
   898 => x"515a5c78",
   899 => x"872484e8",
   900 => x"3862822a",
   901 => x"70810651",
   902 => x"5978802e",
   903 => x"80f83867",
   904 => x"62315a80",
   905 => x"7a2580ee",
   906 => x"38907a25",
   907 => x"b43882b8",
   908 => x"f87c0c90",
   909 => x"0b841d0c",
   910 => x"83b73d08",
   911 => x"900583b8",
   912 => x"3d0c881c",
   913 => x"83b73d08",
   914 => x"811183b9",
   915 => x"3d0c8111",
   916 => x"515a5c78",
   917 => x"87248489",
   918 => x"38f01a5a",
   919 => x"799024ce",
   920 => x"3882b8f8",
   921 => x"7c0c7984",
   922 => x"1d0c83b7",
   923 => x"3d081a83",
   924 => x"b83d0c83",
   925 => x"b63d0881",
   926 => x"1183b83d",
   927 => x"0c811151",
   928 => x"59877925",
   929 => x"913883be",
   930 => x"3ddc0552",
   931 => x"6651f6f9",
   932 => x"3f800884",
   933 => x"89386159",
   934 => x"61682583",
   935 => x"38675968",
   936 => x"194983b7",
   937 => x"3d0883e4",
   938 => x"38800b83",
   939 => x"b73d0c65",
   940 => x"5c69802e",
   941 => x"f88e3869",
   942 => x"5180e8b8",
   943 => x"3f807d5f",
   944 => x"4af88339",
   945 => x"62900743",
   946 => x"62842a70",
   947 => x"81065159",
   948 => x"78939938",
   949 => x"62862a70",
   950 => x"81065159",
   951 => x"78802e93",
   952 => x"8b386465",
   953 => x"84058212",
   954 => x"225d4659",
   955 => x"805f800b",
   956 => x"83be3d34",
   957 => x"facc3962",
   958 => x"90074362",
   959 => x"842a7081",
   960 => x"06515978",
   961 => x"92f43862",
   962 => x"862a7081",
   963 => x"06515978",
   964 => x"802e92e6",
   965 => x"38646584",
   966 => x"05710890",
   967 => x"2b70902c",
   968 => x"515d4659",
   969 => x"807b2489",
   970 => x"a538815f",
   971 => x"fa943964",
   972 => x"65840571",
   973 => x"084a4659",
   974 => x"678025f9",
   975 => x"99386730",
   976 => x"48628407",
   977 => x"7d335b43",
   978 => x"f98f3981",
   979 => x"1d5d6290",
   980 => x"077d335b",
   981 => x"43f98239",
   982 => x"7f802e9e",
   983 => x"ff3882ce",
   984 => x"3d5e7f7e",
   985 => x"34815f80",
   986 => x"0b83be3d",
   987 => x"34fa9a39",
   988 => x"83be3ddc",
   989 => x"05526651",
   990 => x"f58f3f80",
   991 => x"08829f38",
   992 => x"65f01b5b",
   993 => x"5cfae539",
   994 => x"83be3ddc",
   995 => x"05526651",
   996 => x"f4f73f80",
   997 => x"08828738",
   998 => x"65f01b5b",
   999 => x"5cfbfc39",
  1000 => x"6762315a",
  1001 => x"807a25fb",
  1002 => x"b538907a",
  1003 => x"25b43882",
  1004 => x"b9887c0c",
  1005 => x"900b841d",
  1006 => x"0c83b73d",
  1007 => x"08900583",
  1008 => x"b83d0c88",
  1009 => x"1c83b73d",
  1010 => x"08811183",
  1011 => x"b93d0c81",
  1012 => x"11515a5c",
  1013 => x"78872480",
  1014 => x"d138f01a",
  1015 => x"5a799024",
  1016 => x"ce3882b9",
  1017 => x"887c0c79",
  1018 => x"841d0c83",
  1019 => x"b73d081a",
  1020 => x"83b83d0c",
  1021 => x"881c83b7",
  1022 => x"3d088111",
  1023 => x"83b93d0c",
  1024 => x"8111515a",
  1025 => x"5c877925",
  1026 => x"fad43883",
  1027 => x"be3ddc05",
  1028 => x"526651f3",
  1029 => x"f43f8008",
  1030 => x"81843865",
  1031 => x"6460315b",
  1032 => x"5c798024",
  1033 => x"fac238fb",
  1034 => x"b13983be",
  1035 => x"3ddc0552",
  1036 => x"6651f3d5",
  1037 => x"3f800880",
  1038 => x"e53865f0",
  1039 => x"1b5b5cff",
  1040 => x"9c3983be",
  1041 => x"3ddc0552",
  1042 => x"6651f3bd",
  1043 => x"3f800880",
  1044 => x"cd38655c",
  1045 => x"6081802e",
  1046 => x"098106fa",
  1047 => x"8138fec0",
  1048 => x"3983be3d",
  1049 => x"dc055266",
  1050 => x"51f39e3f",
  1051 => x"8008af38",
  1052 => x"65f01b5b",
  1053 => x"5cfbe539",
  1054 => x"83be3ddc",
  1055 => x"05526651",
  1056 => x"f3873f80",
  1057 => x"08983865",
  1058 => x"5cfb8639",
  1059 => x"83be3ddc",
  1060 => x"05526651",
  1061 => x"f2f33f80",
  1062 => x"08802efc",
  1063 => x"8c386980",
  1064 => x"2e873869",
  1065 => x"5180e4cc",
  1066 => x"3f668c05",
  1067 => x"2270862a",
  1068 => x"7081066b",
  1069 => x"5d515a47",
  1070 => x"78802ef5",
  1071 => x"be38ff59",
  1072 => x"f5bb397c",
  1073 => x"337081ff",
  1074 => x"065a5a78",
  1075 => x"80ec2efc",
  1076 => x"fa386290",
  1077 => x"077a81ff",
  1078 => x"06811f5f",
  1079 => x"4143f681",
  1080 => x"397c7081",
  1081 => x"055e3340",
  1082 => x"7faa2e9c",
  1083 => x"cd388060",
  1084 => x"d0057143",
  1085 => x"5a5a7889",
  1086 => x"26f5e638",
  1087 => x"79101010",
  1088 => x"7a100560",
  1089 => x"05d0057d",
  1090 => x"7081055f",
  1091 => x"33d0115b",
  1092 => x"415a8979",
  1093 => x"27e63879",
  1094 => x"4179ff25",
  1095 => x"f5c338ff",
  1096 => x"41f5be39",
  1097 => x"64658405",
  1098 => x"71085d46",
  1099 => x"59820b82",
  1100 => x"bc986472",
  1101 => x"07454f5f",
  1102 => x"80f84080",
  1103 => x"0b83be3d",
  1104 => x"34f5ff39",
  1105 => x"897b27a4",
  1106 => x"38ff1e5e",
  1107 => x"8a527a51",
  1108 => x"81f29d3f",
  1109 => x"8008b005",
  1110 => x"59787e34",
  1111 => x"8a527a51",
  1112 => x"81f1e73f",
  1113 => x"80085b7a",
  1114 => x"8926de38",
  1115 => x"ff1eb01c",
  1116 => x"5a5e787e",
  1117 => x"3483be3d",
  1118 => x"707f31ff",
  1119 => x"9c05405b",
  1120 => x"f68739ff",
  1121 => x"1e7b8f06",
  1122 => x"6f055a5e",
  1123 => x"78337e34",
  1124 => x"7a842a5b",
  1125 => x"7a802edd",
  1126 => x"38ff1e7b",
  1127 => x"8f066f05",
  1128 => x"5a5e7833",
  1129 => x"7e347a84",
  1130 => x"2a5b7ad7",
  1131 => x"38c73962",
  1132 => x"80c0077d",
  1133 => x"335b43f4",
  1134 => x"a03960ff",
  1135 => x"2e99e138",
  1136 => x"7f80e732",
  1137 => x"70307072",
  1138 => x"07802562",
  1139 => x"80c73270",
  1140 => x"30707207",
  1141 => x"80257307",
  1142 => x"53545e51",
  1143 => x"5b597980",
  1144 => x"2e863860",
  1145 => x"83388141",
  1146 => x"64658805",
  1147 => x"84120872",
  1148 => x"087083bf",
  1149 => x"3d0c7183",
  1150 => x"c03d0c54",
  1151 => x"54465981",
  1152 => x"92e63f80",
  1153 => x"08802e91",
  1154 => x"eb388059",
  1155 => x"80795454",
  1156 => x"83ba3d08",
  1157 => x"83bc3d08",
  1158 => x"5b517952",
  1159 => x"81e6e13f",
  1160 => x"800b8008",
  1161 => x"2484d838",
  1162 => x"82bcac5e",
  1163 => x"835ff4d9",
  1164 => x"3982ce3d",
  1165 => x"5e7f80c3",
  1166 => x"2e8f3862",
  1167 => x"842a7081",
  1168 => x"06515978",
  1169 => x"802e82f6",
  1170 => x"38885380",
  1171 => x"52b43d70",
  1172 => x"525980f0",
  1173 => x"883f7854",
  1174 => x"64658405",
  1175 => x"7108557f",
  1176 => x"546c5346",
  1177 => x"599ab83f",
  1178 => x"80085f80",
  1179 => x"08ff2efc",
  1180 => x"ad38800b",
  1181 => x"83be3d34",
  1182 => x"f48f3982",
  1183 => x"bcb06384",
  1184 => x"2a708106",
  1185 => x"515a4e78",
  1186 => x"82893862",
  1187 => x"862a7081",
  1188 => x"06515978",
  1189 => x"802e81fb",
  1190 => x"38646584",
  1191 => x"05821222",
  1192 => x"5d465982",
  1193 => x"6381065a",
  1194 => x"5f7a802e",
  1195 => x"f38e3878",
  1196 => x"802ef388",
  1197 => x"38627f07",
  1198 => x"43800b83",
  1199 => x"be3d34f3",
  1200 => x"8139800b",
  1201 => x"83be3d34",
  1202 => x"64658405",
  1203 => x"71084046",
  1204 => x"597d802e",
  1205 => x"97cf387f",
  1206 => x"80d32e81",
  1207 => x"ff386284",
  1208 => x"2a708106",
  1209 => x"51597881",
  1210 => x"f3388061",
  1211 => x"24f39138",
  1212 => x"60537852",
  1213 => x"7d5180ec",
  1214 => x"823f605f",
  1215 => x"8008802e",
  1216 => x"f3873880",
  1217 => x"087e315f",
  1218 => x"607f25f2",
  1219 => x"fc38605f",
  1220 => x"f2f73962",
  1221 => x"842a7081",
  1222 => x"06515978",
  1223 => x"8d9d3862",
  1224 => x"862a7081",
  1225 => x"06515978",
  1226 => x"802e8d8f",
  1227 => x"38646584",
  1228 => x"05710852",
  1229 => x"46596879",
  1230 => x"237c5eef",
  1231 => x"8939ab0b",
  1232 => x"83be3d34",
  1233 => x"7c335af1",
  1234 => x"9039805a",
  1235 => x"79101010",
  1236 => x"7a100560",
  1237 => x"05d0057d",
  1238 => x"7081055f",
  1239 => x"33d0115b",
  1240 => x"415a8979",
  1241 => x"27e63879",
  1242 => x"48f0f639",
  1243 => x"62818007",
  1244 => x"7d335b43",
  1245 => x"f0e33962",
  1246 => x"88077d33",
  1247 => x"5b43f0d9",
  1248 => x"3982bc98",
  1249 => x"63842a70",
  1250 => x"8106515a",
  1251 => x"4e78802e",
  1252 => x"fdf93864",
  1253 => x"65840571",
  1254 => x"085d4659",
  1255 => x"fe853962",
  1256 => x"81077d33",
  1257 => x"5b43f0b1",
  1258 => x"3983bd3d",
  1259 => x"335978f0",
  1260 => x"a538a00b",
  1261 => x"83be3d34",
  1262 => x"7c335af0",
  1263 => x"9c396465",
  1264 => x"84054659",
  1265 => x"8319337e",
  1266 => x"34815ff7",
  1267 => x"9a397a30",
  1268 => x"5bad0b83",
  1269 => x"be3d3481",
  1270 => x"5ff0e739",
  1271 => x"7da23d0c",
  1272 => x"80705c5f",
  1273 => x"88537e52",
  1274 => x"a63d7052",
  1275 => x"5a80eced",
  1276 => x"3f7e6124",
  1277 => x"8198387a",
  1278 => x"1010a23d",
  1279 => x"08055978",
  1280 => x"08802eaf",
  1281 => x"38795478",
  1282 => x"085383be",
  1283 => x"3dfcc005",
  1284 => x"526a5197",
  1285 => x"8a3f8008",
  1286 => x"ff2ef982",
  1287 => x"3880081f",
  1288 => x"59786124",
  1289 => x"8e38811b",
  1290 => x"79405b78",
  1291 => x"612e0981",
  1292 => x"06c5387e",
  1293 => x"802ef0d1",
  1294 => x"38811f52",
  1295 => x"6a5180dd",
  1296 => x"c43f8008",
  1297 => x"4a800880",
  1298 => x"2ef8de38",
  1299 => x"88538052",
  1300 => x"795180ec",
  1301 => x"883f7955",
  1302 => x"7e5483be",
  1303 => x"3df38c05",
  1304 => x"5369526a",
  1305 => x"5197a03f",
  1306 => x"80087f2e",
  1307 => x"098106f8",
  1308 => x"ad38696a",
  1309 => x"8008055a",
  1310 => x"5e807934",
  1311 => x"f08b39ad",
  1312 => x"0b83be3d",
  1313 => x"3482bcac",
  1314 => x"5e835fef",
  1315 => x"fc397955",
  1316 => x"7e5483be",
  1317 => x"3df38c05",
  1318 => x"537e526a",
  1319 => x"5196e83f",
  1320 => x"80085f80",
  1321 => x"08ff2ef7",
  1322 => x"f5387da2",
  1323 => x"3d0cff83",
  1324 => x"39620a10",
  1325 => x"0a708106",
  1326 => x"51597880",
  1327 => x"2eefe738",
  1328 => x"61820542",
  1329 => x"efe03962",
  1330 => x"0a100a70",
  1331 => x"81065159",
  1332 => x"78802ef1",
  1333 => x"8238b00b",
  1334 => x"82ce3d34",
  1335 => x"7f028405",
  1336 => x"8ab10534",
  1337 => x"83be3dfc",
  1338 => x"bc057c0c",
  1339 => x"820b841d",
  1340 => x"0c83b73d",
  1341 => x"08820583",
  1342 => x"b83d0c88",
  1343 => x"1c83b73d",
  1344 => x"08811183",
  1345 => x"b93d0c81",
  1346 => x"11515a5c",
  1347 => x"877925f0",
  1348 => x"c638f6ae",
  1349 => x"3980e560",
  1350 => x"2582fe38",
  1351 => x"80598079",
  1352 => x"545483ba",
  1353 => x"3d0883bc",
  1354 => x"3d085b51",
  1355 => x"795281db",
  1356 => x"913f8008",
  1357 => x"86d63882",
  1358 => x"bcc47c0c",
  1359 => x"810b841d",
  1360 => x"0c83b73d",
  1361 => x"08810583",
  1362 => x"b83d0c88",
  1363 => x"1c83b73d",
  1364 => x"08811183",
  1365 => x"b93d0c81",
  1366 => x"11515a5c",
  1367 => x"78872481",
  1368 => x"ac38a43d",
  1369 => x"085b7aa6",
  1370 => x"3d08248b",
  1371 => x"38628106",
  1372 => x"5978802e",
  1373 => x"f19b386b",
  1374 => x"7c0c810b",
  1375 => x"841d0c83",
  1376 => x"b73d0881",
  1377 => x"0583b83d",
  1378 => x"0c881c83",
  1379 => x"b73d0881",
  1380 => x"1183b93d",
  1381 => x"0c811151",
  1382 => x"5a5c7887",
  1383 => x"24819b38",
  1384 => x"ff1b5a80",
  1385 => x"7a25f0e9",
  1386 => x"38907a25",
  1387 => x"b43882b9",
  1388 => x"887c0c90",
  1389 => x"0b841d0c",
  1390 => x"83b73d08",
  1391 => x"900583b8",
  1392 => x"3d0c881c",
  1393 => x"83b73d08",
  1394 => x"811183b9",
  1395 => x"3d0c8111",
  1396 => x"515a5c78",
  1397 => x"872480ca",
  1398 => x"38f01a5a",
  1399 => x"799024ce",
  1400 => x"3882b988",
  1401 => x"7c0c7984",
  1402 => x"1d0c83b7",
  1403 => x"3d081a83",
  1404 => x"b83d0c88",
  1405 => x"1c83b73d",
  1406 => x"08811183",
  1407 => x"b93d0c81",
  1408 => x"11515a5c",
  1409 => x"877925f0",
  1410 => x"8838f4ec",
  1411 => x"3983be3d",
  1412 => x"dc055266",
  1413 => x"51e7f23f",
  1414 => x"8008f582",
  1415 => x"38655cfe",
  1416 => x"c13983be",
  1417 => x"3ddc0552",
  1418 => x"6651e7dd",
  1419 => x"3f8008f4",
  1420 => x"ed3865f0",
  1421 => x"1b5b5cff",
  1422 => x"a33983be",
  1423 => x"3ddc0552",
  1424 => x"6651e7c5",
  1425 => x"3f8008f4",
  1426 => x"d53865a5",
  1427 => x"3d08ff05",
  1428 => x"5b5c7980",
  1429 => x"24fed238",
  1430 => x"efb73983",
  1431 => x"be3ddc05",
  1432 => x"526651e7",
  1433 => x"a43f8008",
  1434 => x"f4b43865",
  1435 => x"83be3d33",
  1436 => x"5c5cedab",
  1437 => x"397ef5fd",
  1438 => x"38628106",
  1439 => x"5978802e",
  1440 => x"f5f33802",
  1441 => x"8d8f055e",
  1442 => x"b07e3483",
  1443 => x"be3d707f",
  1444 => x"31ff9c05",
  1445 => x"405bebf1",
  1446 => x"39a43d08",
  1447 => x"5b817b25",
  1448 => x"8382387d",
  1449 => x"7081055f",
  1450 => x"3382ce3d",
  1451 => x"34ae0284",
  1452 => x"058ab105",
  1453 => x"3483be3d",
  1454 => x"fcbc057c",
  1455 => x"0c820b84",
  1456 => x"1d0c83b7",
  1457 => x"3d088205",
  1458 => x"83b83d0c",
  1459 => x"881c83b7",
  1460 => x"3d088111",
  1461 => x"83b93d0c",
  1462 => x"8111515a",
  1463 => x"5c788724",
  1464 => x"80fd3880",
  1465 => x"59807954",
  1466 => x"5483ba3d",
  1467 => x"0883bc3d",
  1468 => x"085b5179",
  1469 => x"5281d9b4",
  1470 => x"3f800880",
  1471 => x"2e819138",
  1472 => x"7d7c0cff",
  1473 => x"1b841d0c",
  1474 => x"83b73d08",
  1475 => x"1bff0583",
  1476 => x"b83d0c88",
  1477 => x"1c83b73d",
  1478 => x"08811183",
  1479 => x"b93d0c81",
  1480 => x"11515a5c",
  1481 => x"78872481",
  1482 => x"d13883be",
  1483 => x"3de8057c",
  1484 => x"0c6c841d",
  1485 => x"0c83b73d",
  1486 => x"086d0583",
  1487 => x"b83d0c88",
  1488 => x"1c83b73d",
  1489 => x"08811183",
  1490 => x"b93d0c81",
  1491 => x"11515a5c",
  1492 => x"877925ed",
  1493 => x"bc3883be",
  1494 => x"3ddc0552",
  1495 => x"f2a03983",
  1496 => x"be3ddc05",
  1497 => x"526651e5",
  1498 => x"a03f8008",
  1499 => x"f2b03865",
  1500 => x"a53d085c",
  1501 => x"5c805980",
  1502 => x"79545483",
  1503 => x"ba3d0883",
  1504 => x"bc3d085b",
  1505 => x"51795281",
  1506 => x"d8a23f80",
  1507 => x"08fef138",
  1508 => x"ff1b5a80",
  1509 => x"7a25ff92",
  1510 => x"38907a25",
  1511 => x"b43882b9",
  1512 => x"887c0c90",
  1513 => x"0b841d0c",
  1514 => x"83b73d08",
  1515 => x"900583b8",
  1516 => x"3d0c881c",
  1517 => x"83b73d08",
  1518 => x"811183b9",
  1519 => x"3d0c8111",
  1520 => x"515a5c78",
  1521 => x"872483db",
  1522 => x"38f01a5a",
  1523 => x"799024ce",
  1524 => x"3882b988",
  1525 => x"7c0c7984",
  1526 => x"1d0c83b7",
  1527 => x"3d081a83",
  1528 => x"b83d0c88",
  1529 => x"1c83b73d",
  1530 => x"08811183",
  1531 => x"b93d0c81",
  1532 => x"11515a5c",
  1533 => x"877925fe",
  1534 => x"b13883be",
  1535 => x"3ddc0552",
  1536 => x"6651e485",
  1537 => x"3f8008f1",
  1538 => x"95386583",
  1539 => x"bf3de805",
  1540 => x"710c6d84",
  1541 => x"120c83b8",
  1542 => x"3d086e05",
  1543 => x"83b93d0c",
  1544 => x"5cfe9c39",
  1545 => x"62810659",
  1546 => x"78fcf838",
  1547 => x"7d7c0c81",
  1548 => x"0b841d0c",
  1549 => x"83b73d08",
  1550 => x"810583b8",
  1551 => x"3d0c881c",
  1552 => x"83b73d08",
  1553 => x"811183b9",
  1554 => x"3d0c8111",
  1555 => x"515a5c87",
  1556 => x"7925fdd6",
  1557 => x"3883be3d",
  1558 => x"dc0552ff",
  1559 => x"a3396465",
  1560 => x"84057108",
  1561 => x"5d465981",
  1562 => x"5fe7d139",
  1563 => x"64658405",
  1564 => x"71085d46",
  1565 => x"59805fec",
  1566 => x"f5396465",
  1567 => x"84057108",
  1568 => x"5d46597a",
  1569 => x"8025eda2",
  1570 => x"38f6c339",
  1571 => x"a53d085a",
  1572 => x"807a2589",
  1573 => x"c638a43d",
  1574 => x"085b7a7a",
  1575 => x"2482dd38",
  1576 => x"7d7c0c7a",
  1577 => x"841d0c83",
  1578 => x"b73d081b",
  1579 => x"83b83d0c",
  1580 => x"881c83b7",
  1581 => x"3d088111",
  1582 => x"83b93d0c",
  1583 => x"8111515a",
  1584 => x"5c788724",
  1585 => x"81b63879",
  1586 => x"7b315a80",
  1587 => x"7a2580f3",
  1588 => x"38907a25",
  1589 => x"b43882b9",
  1590 => x"887c0c90",
  1591 => x"0b841d0c",
  1592 => x"83b73d08",
  1593 => x"900583b8",
  1594 => x"3d0c881c",
  1595 => x"83b73d08",
  1596 => x"811183b9",
  1597 => x"3d0c8111",
  1598 => x"515a5c78",
  1599 => x"872480e4",
  1600 => x"38f01a5a",
  1601 => x"799024ce",
  1602 => x"3882b988",
  1603 => x"7c0c7984",
  1604 => x"1d0c83b7",
  1605 => x"3d081a83",
  1606 => x"b83d0c88",
  1607 => x"1c83b73d",
  1608 => x"08811183",
  1609 => x"b93d0c81",
  1610 => x"11515a5c",
  1611 => x"87792593",
  1612 => x"3883be3d",
  1613 => x"dc055266",
  1614 => x"51e1ce3f",
  1615 => x"8008eede",
  1616 => x"38655c62",
  1617 => x"81065978",
  1618 => x"802ee9c5",
  1619 => x"3882bcc8",
  1620 => x"7c0c810b",
  1621 => x"841d0c83",
  1622 => x"b73d0881",
  1623 => x"0583b83d",
  1624 => x"0cfbdc39",
  1625 => x"83be3ddc",
  1626 => x"05526651",
  1627 => x"e19b3f80",
  1628 => x"08eeab38",
  1629 => x"65f01b5b",
  1630 => x"5cff8939",
  1631 => x"83be3ddc",
  1632 => x"05526651",
  1633 => x"e1833f80",
  1634 => x"08ee9338",
  1635 => x"65a63d08",
  1636 => x"a63d0871",
  1637 => x"7131525d",
  1638 => x"5b5c7980",
  1639 => x"24feb238",
  1640 => x"ffa13983",
  1641 => x"be3ddc05",
  1642 => x"526651e0",
  1643 => x"dc3f8008",
  1644 => x"edec3865",
  1645 => x"f01b5b5c",
  1646 => x"fc923964",
  1647 => x"65840571",
  1648 => x"086b710c",
  1649 => x"527e4046",
  1650 => x"59e1fb39",
  1651 => x"7ee5ad38",
  1652 => x"ff1e7bb7",
  1653 => x"06b0075b",
  1654 => x"5e797e34",
  1655 => x"7a832a5b",
  1656 => x"7aee3862",
  1657 => x"81065978",
  1658 => x"802eef89",
  1659 => x"3879b02e",
  1660 => x"ef8338ff",
  1661 => x"1e5eb07e",
  1662 => x"34f99039",
  1663 => x"7d7c0c79",
  1664 => x"841d0c83",
  1665 => x"b73d081a",
  1666 => x"83b83d0c",
  1667 => x"881c83b7",
  1668 => x"3d088111",
  1669 => x"83b93d0c",
  1670 => x"8111515a",
  1671 => x"5c788724",
  1672 => x"818b3879",
  1673 => x"1e82bcc8",
  1674 => x"7d0c5e81",
  1675 => x"0b841d0c",
  1676 => x"83b73d08",
  1677 => x"810583b8",
  1678 => x"3d0c881c",
  1679 => x"83b73d08",
  1680 => x"811183b9",
  1681 => x"3d0c8111",
  1682 => x"515a5c78",
  1683 => x"8724b038",
  1684 => x"7d7c0ca4",
  1685 => x"3d087a31",
  1686 => x"70841e0c",
  1687 => x"83b83d08",
  1688 => x"0583b83d",
  1689 => x"0c881c83",
  1690 => x"b73d0881",
  1691 => x"1183b93d",
  1692 => x"0c811151",
  1693 => x"5a5c8779",
  1694 => x"25e79638",
  1695 => x"ebfa3983",
  1696 => x"be3ddc05",
  1697 => x"526651df",
  1698 => x"803f8008",
  1699 => x"ec903865",
  1700 => x"a63d087f",
  1701 => x"720ca63d",
  1702 => x"08713170",
  1703 => x"84140c83",
  1704 => x"ba3d0805",
  1705 => x"83ba3d0c",
  1706 => x"5b5cffb9",
  1707 => x"3983be3d",
  1708 => x"dc055266",
  1709 => x"51ded23f",
  1710 => x"8008ebe2",
  1711 => x"3865a63d",
  1712 => x"087f1182",
  1713 => x"bcc8730c",
  1714 => x"405b5c81",
  1715 => x"0b841d0c",
  1716 => x"83b73d08",
  1717 => x"810583b8",
  1718 => x"3d0c881c",
  1719 => x"83b73d08",
  1720 => x"811183b9",
  1721 => x"3d0c8111",
  1722 => x"515a5c87",
  1723 => x"7925fee0",
  1724 => x"38ff8c39",
  1725 => x"83ba3d08",
  1726 => x"83bc3d08",
  1727 => x"5b517952",
  1728 => x"8181963f",
  1729 => x"82bccc5e",
  1730 => x"835f8008",
  1731 => x"e2fb3862",
  1732 => x"82800783",
  1733 => x"bb3d0883",
  1734 => x"bd3d0863",
  1735 => x"83c03daa",
  1736 => x"3da53d0c",
  1737 => x"5f45415f",
  1738 => x"43830ba1",
  1739 => x"3d0c7f80",
  1740 => x"e62ea738",
  1741 => x"80085a7f",
  1742 => x"80e52e83",
  1743 => x"a7388008",
  1744 => x"597f80c5",
  1745 => x"2e83ad38",
  1746 => x"79790759",
  1747 => x"78802e85",
  1748 => x"38608105",
  1749 => x"42820ba1",
  1750 => x"3d0c7db3",
  1751 => x"3d0c7eb4",
  1752 => x"3d0c800b",
  1753 => x"b33d0824",
  1754 => x"879a3880",
  1755 => x"7b3483be",
  1756 => x"3df39411",
  1757 => x"59f39005",
  1758 => x"576e5661",
  1759 => x"556f547d",
  1760 => x"527e536a",
  1761 => x"5196cf3f",
  1762 => x"80086080",
  1763 => x"e7327030",
  1764 => x"7072079f",
  1765 => x"2a515b5b",
  1766 => x"a13d0c7f",
  1767 => x"80c72e85",
  1768 => x"387881ce",
  1769 => x"38628106",
  1770 => x"597881c6",
  1771 => x"38a33d08",
  1772 => x"5978a13d",
  1773 => x"0831a53d",
  1774 => x"0c6f6080",
  1775 => x"e7327030",
  1776 => x"70720780",
  1777 => x"256380c7",
  1778 => x"32703070",
  1779 => x"72078025",
  1780 => x"73075354",
  1781 => x"5f515c5a",
  1782 => x"5e79802e",
  1783 => x"85d038a5",
  1784 => x"3d085afc",
  1785 => x"7a258738",
  1786 => x"607a2582",
  1787 => x"9d3880e5",
  1788 => x"597f80e7",
  1789 => x"2e843880",
  1790 => x"c5597840",
  1791 => x"7f80e524",
  1792 => x"85b338ff",
  1793 => x"1a70a73d",
  1794 => x"0c83b93d",
  1795 => x"715d435a",
  1796 => x"7f623402",
  1797 => x"8ddd055f",
  1798 => x"807a2486",
  1799 => x"8438ab7f",
  1800 => x"34028dde",
  1801 => x"05b33d70",
  1802 => x"5c425f89",
  1803 => x"7b2580fb",
  1804 => x"38ff1a5a",
  1805 => x"8a527a51",
  1806 => x"d6d73f80",
  1807 => x"08b00559",
  1808 => x"787a348a",
  1809 => x"527a51d5",
  1810 => x"963f8008",
  1811 => x"5b800889",
  1812 => x"24df38ff",
  1813 => x"1a8008b0",
  1814 => x"055a5a78",
  1815 => x"7a347961",
  1816 => x"2780d938",
  1817 => x"79708105",
  1818 => x"5b337f70",
  1819 => x"81054134",
  1820 => x"ed398008",
  1821 => x"62055b7f",
  1822 => x"80e62e80",
  1823 => x"fc388059",
  1824 => x"80795454",
  1825 => x"7d517e52",
  1826 => x"81ccb73f",
  1827 => x"80088538",
  1828 => x"7aa43d0c",
  1829 => x"a33d0859",
  1830 => x"787b27fe",
  1831 => x"9438b079",
  1832 => x"34a33d08",
  1833 => x"8105a43d",
  1834 => x"0cea39b0",
  1835 => x"7f708105",
  1836 => x"4134b01b",
  1837 => x"59787f70",
  1838 => x"81054134",
  1839 => x"7e6231a5",
  1840 => x"3d087012",
  1841 => x"415a4d81",
  1842 => x"792580ff",
  1843 => x"38811f5f",
  1844 => x"83bc3d33",
  1845 => x"5978802e",
  1846 => x"dfaf38ad",
  1847 => x"0b83be3d",
  1848 => x"34dfa639",
  1849 => x"810b8008",
  1850 => x"5a5a7f80",
  1851 => x"c52e0981",
  1852 => x"06fcd538",
  1853 => x"8159fcd0",
  1854 => x"39800833",
  1855 => x"5978b02e",
  1856 => x"a8386e08",
  1857 => x"7b055bfe",
  1858 => x"f53980e7",
  1859 => x"40a43d08",
  1860 => x"59787a24",
  1861 => x"83f93879",
  1862 => x"6381065a",
  1863 => x"5f78802e",
  1864 => x"ffae3881",
  1865 => x"1a5fffa8",
  1866 => x"39805980",
  1867 => x"7954547d",
  1868 => x"517e5281",
  1869 => x"ccf63f80",
  1870 => x"08802ec6",
  1871 => x"38816231",
  1872 => x"70a13d08",
  1873 => x"0c7b055b",
  1874 => x"feb43962",
  1875 => x"81065978",
  1876 => x"802efefc",
  1877 => x"38811f5f",
  1878 => x"fef63982",
  1879 => x"bcc47c0c",
  1880 => x"810b841d",
  1881 => x"0c83b73d",
  1882 => x"08810583",
  1883 => x"b83d0c88",
  1884 => x"1c83b73d",
  1885 => x"08811183",
  1886 => x"b93d0c81",
  1887 => x"11515a5c",
  1888 => x"78872481",
  1889 => x"e0387989",
  1890 => x"38a43d08",
  1891 => x"802ee181",
  1892 => x"386b7c0c",
  1893 => x"810b841d",
  1894 => x"0c83b73d",
  1895 => x"08810583",
  1896 => x"b83d0c88",
  1897 => x"1c83b73d",
  1898 => x"08811183",
  1899 => x"b93d0c81",
  1900 => x"11515a5c",
  1901 => x"78872481",
  1902 => x"c5387930",
  1903 => x"5a807a25",
  1904 => x"80f33890",
  1905 => x"7a25b438",
  1906 => x"82b9887c",
  1907 => x"0c900b84",
  1908 => x"1d0c83b7",
  1909 => x"3d089005",
  1910 => x"83b83d0c",
  1911 => x"881c83b7",
  1912 => x"3d088111",
  1913 => x"83b93d0c",
  1914 => x"8111515a",
  1915 => x"5c788724",
  1916 => x"80db38f0",
  1917 => x"1a5a7990",
  1918 => x"24ce3882",
  1919 => x"b9887c0c",
  1920 => x"79841d0c",
  1921 => x"83b73d08",
  1922 => x"1a83b83d",
  1923 => x"0c881c83",
  1924 => x"b73d0881",
  1925 => x"1183b93d",
  1926 => x"0c811151",
  1927 => x"5a5c8779",
  1928 => x"25933883",
  1929 => x"be3ddc05",
  1930 => x"526651d7",
  1931 => x"dc3f8008",
  1932 => x"e4ec3865",
  1933 => x"5c7d7c0c",
  1934 => x"a43d0884",
  1935 => x"1d0c83b7",
  1936 => x"3d08a53d",
  1937 => x"080583b8",
  1938 => x"3d0cf1f3",
  1939 => x"3983be3d",
  1940 => x"dc055266",
  1941 => x"51d7b23f",
  1942 => x"8008e4c2",
  1943 => x"3865f01b",
  1944 => x"5b5cff92",
  1945 => x"3983be3d",
  1946 => x"dc055266",
  1947 => x"51d79a3f",
  1948 => x"8008e4aa",
  1949 => x"3865a63d",
  1950 => x"085b5cfe",
  1951 => x"893983be",
  1952 => x"3ddc0552",
  1953 => x"6651d781",
  1954 => x"3f8008e4",
  1955 => x"913865a6",
  1956 => x"3d087030",
  1957 => x"515b5c79",
  1958 => x"8024fea7",
  1959 => x"38ff9639",
  1960 => x"8641e6c4",
  1961 => x"3982bcd0",
  1962 => x"5e865fdb",
  1963 => x"dc39a53d",
  1964 => x"085afac8",
  1965 => x"397f80e6",
  1966 => x"2e098106",
  1967 => x"fccf3880",
  1968 => x"7a25818d",
  1969 => x"38795f60",
  1970 => x"8b386281",
  1971 => x"06597880",
  1972 => x"2efbfd38",
  1973 => x"601a8105",
  1974 => x"5ffbf539",
  1975 => x"83b73d08",
  1976 => x"8a38800b",
  1977 => x"83b73d0c",
  1978 => x"e3b43983",
  1979 => x"be3ddc05",
  1980 => x"526651d6",
  1981 => x"943f8008",
  1982 => x"e3a43880",
  1983 => x"0b83b73d",
  1984 => x"0ce39b39",
  1985 => x"7d810a32",
  1986 => x"5ead7b34",
  1987 => x"f8e03978",
  1988 => x"7a318205",
  1989 => x"5f807a25",
  1990 => x"fbb63881",
  1991 => x"195ffbb0",
  1992 => x"3979305b",
  1993 => x"ad7f3402",
  1994 => x"8dde05b3",
  1995 => x"3d705c42",
  1996 => x"5f897b25",
  1997 => x"faf538f9",
  1998 => x"f8396465",
  1999 => x"84057108",
  2000 => x"43465960",
  2001 => x"8025d98e",
  2002 => x"38ff7d33",
  2003 => x"5b41d989",
  2004 => x"39608d38",
  2005 => x"62810659",
  2006 => x"815f7880",
  2007 => x"2efaf138",
  2008 => x"6082055f",
  2009 => x"faea39fc",
  2010 => x"3d0d82c0",
  2011 => x"c00855b8",
  2012 => x"1508802e",
  2013 => x"93387854",
  2014 => x"77537652",
  2015 => x"82c0c008",
  2016 => x"51d5b73f",
  2017 => x"863d0d04",
  2018 => x"7451b3fb",
  2019 => x"3f785477",
  2020 => x"53765282",
  2021 => x"c0c00851",
  2022 => x"d5a03f86",
  2023 => x"3d0d04f6",
  2024 => x"3d0d7c7e",
  2025 => x"61595658",
  2026 => x"80567476",
  2027 => x"2e9c3876",
  2028 => x"547e5374",
  2029 => x"52775182",
  2030 => x"b73f8008",
  2031 => x"558008ff",
  2032 => x"2ea23874",
  2033 => x"800c8c3d",
  2034 => x"0d047654",
  2035 => x"75538c3d",
  2036 => x"f4055277",
  2037 => x"5182993f",
  2038 => x"80085580",
  2039 => x"08ff2e09",
  2040 => x"8106e038",
  2041 => x"80770c81",
  2042 => x"8a780c74",
  2043 => x"800c8c3d",
  2044 => x"0d04fd3d",
  2045 => x"0d775476",
  2046 => x"53755282",
  2047 => x"c0c00851",
  2048 => x"ff9d3f85",
  2049 => x"3d0d04ec",
  2050 => x"3d0d6668",
  2051 => x"6a6c6e73",
  2052 => x"5c405d42",
  2053 => x"42426080",
  2054 => x"2e818c38",
  2055 => x"8060085a",
  2056 => x"5d7c7a27",
  2057 => x"80f83893",
  2058 => x"3d5b7b08",
  2059 => x"841d087d",
  2060 => x"567a0855",
  2061 => x"7c546353",
  2062 => x"405efee3",
  2063 => x"3f800858",
  2064 => x"8008ff2e",
  2065 => x"80f13880",
  2066 => x"7a800831",
  2067 => x"56567c75",
  2068 => x"26833881",
  2069 => x"5680087a",
  2070 => x"2780d138",
  2071 => x"75802e80",
  2072 => x"cb388008",
  2073 => x"1d5d6080",
  2074 => x"2ea23880",
  2075 => x"56758008",
  2076 => x"25943875",
  2077 => x"1b557433",
  2078 => x"77708105",
  2079 => x"59348116",
  2080 => x"56777624",
  2081 => x"ee387f08",
  2082 => x"8405600c",
  2083 => x"78708405",
  2084 => x"5a085574",
  2085 => x"802eaf38",
  2086 => x"797d26ff",
  2087 => x"8d387c55",
  2088 => x"74800c96",
  2089 => x"3d0d04ff",
  2090 => x"5afef139",
  2091 => x"7d7c0c7e",
  2092 => x"841d0c7c",
  2093 => x"55ea3981",
  2094 => x"8a620c80",
  2095 => x"7c0c8008",
  2096 => x"800c963d",
  2097 => x"0d046080",
  2098 => x"2e843874",
  2099 => x"600c747c",
  2100 => x"0cff1d80",
  2101 => x"0c963d0d",
  2102 => x"04fc3d0d",
  2103 => x"79557854",
  2104 => x"77537652",
  2105 => x"82c0c008",
  2106 => x"51fe9c3f",
  2107 => x"863d0d04",
  2108 => x"f83d0d7b",
  2109 => x"7d7f82c7",
  2110 => x"c0545957",
  2111 => x"5580f98a",
  2112 => x"3f800881",
  2113 => x"26943874",
  2114 => x"5474802e",
  2115 => x"86387575",
  2116 => x"34815473",
  2117 => x"800c8a3d",
  2118 => x"0d0482bc",
  2119 => x"d85282c7",
  2120 => x"c05180f7",
  2121 => x"d03f8008",
  2122 => x"81c13880",
  2123 => x"08547480",
  2124 => x"2ee13880",
  2125 => x"ff7625d6",
  2126 => x"38ff8016",
  2127 => x"538eff73",
  2128 => x"2784ef38",
  2129 => x"f0801653",
  2130 => x"83efff73",
  2131 => x"2782a938",
  2132 => x"fc808016",
  2133 => x"5380fbff",
  2134 => x"ff732784",
  2135 => x"f7388fff",
  2136 => x"0a1653f7",
  2137 => x"c00a7327",
  2138 => x"85b838ff",
  2139 => x"54c00a76",
  2140 => x"25ffa038",
  2141 => x"75820a06",
  2142 => x"709e2c70",
  2143 => x"fc075151",
  2144 => x"53727570",
  2145 => x"81055734",
  2146 => x"7581fc0a",
  2147 => x"0670982a",
  2148 => x"ff800751",
  2149 => x"53727570",
  2150 => x"81055734",
  2151 => x"7587f080",
  2152 => x"80067092",
  2153 => x"2aff8007",
  2154 => x"51537275",
  2155 => x"70810557",
  2156 => x"34758fe0",
  2157 => x"8006708c",
  2158 => x"2aff8007",
  2159 => x"51537275",
  2160 => x"70810557",
  2161 => x"34759fc0",
  2162 => x"0670862a",
  2163 => x"ff800751",
  2164 => x"53727570",
  2165 => x"81055734",
  2166 => x"75ffbf06",
  2167 => x"ff800753",
  2168 => x"72753486",
  2169 => x"0b800c8a",
  2170 => x"3d0d0482",
  2171 => x"bce05282",
  2172 => x"c7c05180",
  2173 => x"f5ff3f80",
  2174 => x"0881d738",
  2175 => x"7581ff06",
  2176 => x"76882c70",
  2177 => x"81ff0680",
  2178 => x"08575954",
  2179 => x"5874802e",
  2180 => x"fe813876",
  2181 => x"802efdef",
  2182 => x"38800880",
  2183 => x"ff187081",
  2184 => x"ff065154",
  2185 => x"56729e26",
  2186 => x"83388156",
  2187 => x"8008a018",
  2188 => x"7081ff06",
  2189 => x"51545472",
  2190 => x"8f268338",
  2191 => x"81547574",
  2192 => x"07537280",
  2193 => x"2eaa3880",
  2194 => x"08c01954",
  2195 => x"5672be26",
  2196 => x"83388156",
  2197 => x"8008ff80",
  2198 => x"197081ff",
  2199 => x"06515454",
  2200 => x"7280fc26",
  2201 => x"83388154",
  2202 => x"75740753",
  2203 => x"7280d038",
  2204 => x"ff0b800c",
  2205 => x"8a3d0d04",
  2206 => x"fcd08016",
  2207 => x"53ff548f",
  2208 => x"ff7327fd",
  2209 => x"8e387583",
  2210 => x"e0800670",
  2211 => x"8c2ae007",
  2212 => x"51537275",
  2213 => x"70810557",
  2214 => x"34759fc0",
  2215 => x"0670862a",
  2216 => x"ff800751",
  2217 => x"53727570",
  2218 => x"81055734",
  2219 => x"75ffbf06",
  2220 => x"ff800753",
  2221 => x"72753483",
  2222 => x"0b800c8a",
  2223 => x"3d0d0476",
  2224 => x"75708105",
  2225 => x"57347775",
  2226 => x"34825473",
  2227 => x"800c8a3d",
  2228 => x"0d0482bc",
  2229 => x"e85282c7",
  2230 => x"c05180f4",
  2231 => x"983f8008",
  2232 => x"80db3875",
  2233 => x"81ff0676",
  2234 => x"882c7081",
  2235 => x"ff068008",
  2236 => x"57595458",
  2237 => x"74802efc",
  2238 => x"9a387680",
  2239 => x"2efc8838",
  2240 => x"80085381",
  2241 => x"a0772783",
  2242 => x"38815376",
  2243 => x"81ff2efe",
  2244 => x"df388170",
  2245 => x"74065454",
  2246 => x"72802efe",
  2247 => x"d3388008",
  2248 => x"5381a078",
  2249 => x"27833873",
  2250 => x"537781ff",
  2251 => x"2efec138",
  2252 => x"72740653",
  2253 => x"72802efe",
  2254 => x"b738ff83",
  2255 => x"3982bcf0",
  2256 => x"5282c7c0",
  2257 => x"5180f3ad",
  2258 => x"3f8008fb",
  2259 => x"ba388008",
  2260 => x"7681ff06",
  2261 => x"77882c70",
  2262 => x"81ff0659",
  2263 => x"55595981",
  2264 => x"5474802e",
  2265 => x"fbad3875",
  2266 => x"802e8298",
  2267 => x"38df1653",
  2268 => x"7280dd26",
  2269 => x"fdfa38df",
  2270 => x"18537280",
  2271 => x"dd26fdf0",
  2272 => x"3876089c",
  2273 => x"3873770c",
  2274 => x"9b757081",
  2275 => x"055734a4",
  2276 => x"75708105",
  2277 => x"573480c2",
  2278 => x"75708105",
  2279 => x"57348359",
  2280 => x"75757081",
  2281 => x"05573477",
  2282 => x"75348219",
  2283 => x"800c8a3d",
  2284 => x"0d04758f",
  2285 => x"c0067086",
  2286 => x"2ac00751",
  2287 => x"53727570",
  2288 => x"81055734",
  2289 => x"75ffbf06",
  2290 => x"ff800753",
  2291 => x"72753482",
  2292 => x"54fdf839",
  2293 => x"7580f080",
  2294 => x"80067092",
  2295 => x"2af00751",
  2296 => x"53727570",
  2297 => x"81055734",
  2298 => x"758fe080",
  2299 => x"06708c2a",
  2300 => x"ff800751",
  2301 => x"53727570",
  2302 => x"81055734",
  2303 => x"759fc006",
  2304 => x"70862aff",
  2305 => x"80075153",
  2306 => x"72757081",
  2307 => x"05573475",
  2308 => x"ffbf06ff",
  2309 => x"80075372",
  2310 => x"7534840b",
  2311 => x"800c8a3d",
  2312 => x"0d047581",
  2313 => x"c00a0670",
  2314 => x"982af807",
  2315 => x"51537275",
  2316 => x"70810557",
  2317 => x"347587f0",
  2318 => x"80800670",
  2319 => x"922aff80",
  2320 => x"07515372",
  2321 => x"75708105",
  2322 => x"5734758f",
  2323 => x"e0800670",
  2324 => x"8c2aff80",
  2325 => x"07515372",
  2326 => x"75708105",
  2327 => x"5734759f",
  2328 => x"c0067086",
  2329 => x"2aff8007",
  2330 => x"51537275",
  2331 => x"70810557",
  2332 => x"3475ffbf",
  2333 => x"06ff8007",
  2334 => x"53727534",
  2335 => x"850b800c",
  2336 => x"8a3d0d04",
  2337 => x"7608802e",
  2338 => x"9d388008",
  2339 => x"770c9b75",
  2340 => x"70810557",
  2341 => x"34a87570",
  2342 => x"81055734",
  2343 => x"80c27570",
  2344 => x"81055734",
  2345 => x"83597775",
  2346 => x"34811980",
  2347 => x"0c8a3d0d",
  2348 => x"04fa3d0d",
  2349 => x"7882c0c0",
  2350 => x"085455b8",
  2351 => x"1308802e",
  2352 => x"81b6388c",
  2353 => x"15227083",
  2354 => x"ffff0670",
  2355 => x"832a8132",
  2356 => x"70810651",
  2357 => x"55555672",
  2358 => x"802e80dc",
  2359 => x"3873842a",
  2360 => x"81328106",
  2361 => x"57ff5376",
  2362 => x"80f73873",
  2363 => x"822a7081",
  2364 => x"06515372",
  2365 => x"802eb938",
  2366 => x"b0150854",
  2367 => x"73802e9c",
  2368 => x"3880c015",
  2369 => x"5373732e",
  2370 => x"8f387352",
  2371 => x"82c0c008",
  2372 => x"51acde3f",
  2373 => x"8c152256",
  2374 => x"76b0160c",
  2375 => x"75db0653",
  2376 => x"728c1623",
  2377 => x"800b8416",
  2378 => x"0c901508",
  2379 => x"750c7256",
  2380 => x"75880753",
  2381 => x"728c1623",
  2382 => x"90150880",
  2383 => x"2e80c138",
  2384 => x"8c152270",
  2385 => x"81065553",
  2386 => x"739e3872",
  2387 => x"0a100a70",
  2388 => x"81065153",
  2389 => x"72853894",
  2390 => x"15085473",
  2391 => x"88160c80",
  2392 => x"5372800c",
  2393 => x"883d0d04",
  2394 => x"800b8816",
  2395 => x"0c941508",
  2396 => x"3098160c",
  2397 => x"8053ea39",
  2398 => x"7251a88b",
  2399 => x"3ffec439",
  2400 => x"7451b8dc",
  2401 => x"3f8c1522",
  2402 => x"70810655",
  2403 => x"5373802e",
  2404 => x"ffb938d4",
  2405 => x"39ef3d0d",
  2406 => x"63659011",
  2407 => x"085e4040",
  2408 => x"80537b60",
  2409 => x"90050824",
  2410 => x"81b33894",
  2411 => x"1f70ff1e",
  2412 => x"70822b73",
  2413 => x"11649405",
  2414 => x"705c435f",
  2415 => x"61057008",
  2416 => x"7f088105",
  2417 => x"57555c5e",
  2418 => x"425781c8",
  2419 => x"fd3f8008",
  2420 => x"5d800881",
  2421 => x"8f387e52",
  2422 => x"7f5180d5",
  2423 => x"f53f800b",
  2424 => x"80082480",
  2425 => x"f638811d",
  2426 => x"5d80707f",
  2427 => x"635a585b",
  2428 => x"58767084",
  2429 => x"05580870",
  2430 => x"83ffff06",
  2431 => x"7b057190",
  2432 => x"2a71902a",
  2433 => x"0570902a",
  2434 => x"5d5283ff",
  2435 => x"ff068218",
  2436 => x"22707231",
  2437 => x"1b585b54",
  2438 => x"83ffff06",
  2439 => x"76227072",
  2440 => x"3177902c",
  2441 => x"0570902c",
  2442 => x"5b524353",
  2443 => x"72762374",
  2444 => x"82172384",
  2445 => x"16567a77",
  2446 => x"27ffb638",
  2447 => x"7b10101e",
  2448 => x"59780897",
  2449 => x"38fc1959",
  2450 => x"7d79278a",
  2451 => x"38780886",
  2452 => x"38ff1c5c",
  2453 => x"f0397b60",
  2454 => x"90050c7c",
  2455 => x"5372800c",
  2456 => x"933d0d04",
  2457 => x"80705b58",
  2458 => x"76708405",
  2459 => x"58087083",
  2460 => x"ffff0670",
  2461 => x"7f291c72",
  2462 => x"902a6029",
  2463 => x"71902a05",
  2464 => x"70902a5e",
  2465 => x"5283ffff",
  2466 => x"06821922",
  2467 => x"7072311c",
  2468 => x"59455283",
  2469 => x"ffff0677",
  2470 => x"22707231",
  2471 => x"78902c05",
  2472 => x"70902c5c",
  2473 => x"52565153",
  2474 => x"72762374",
  2475 => x"82172384",
  2476 => x"16567a77",
  2477 => x"27ffb138",
  2478 => x"7808fe9a",
  2479 => x"38fc1959",
  2480 => x"7d79278a",
  2481 => x"38780886",
  2482 => x"38ff1c5c",
  2483 => x"f0397b60",
  2484 => x"90050cfe",
  2485 => x"81398c08",
  2486 => x"c83d0dbc",
  2487 => x"3d0880c0",
  2488 => x"3d0880c2",
  2489 => x"3d0880c5",
  2490 => x"3d0880c7",
  2491 => x"3d088c0c",
  2492 => x"5d4b4340",
  2493 => x"800bbe3d",
  2494 => x"0880c03d",
  2495 => x"085bba3d",
  2496 => x"0c79bb3d",
  2497 => x"0c6080c0",
  2498 => x"05085748",
  2499 => x"75682e09",
  2500 => x"810680d9",
  2501 => x"38b83d08",
  2502 => x"57807724",
  2503 => x"80f93867",
  2504 => x"7a0c769f",
  2505 => x"fe0a0656",
  2506 => x"759ffe0a",
  2507 => x"2e818538",
  2508 => x"b83d08ba",
  2509 => x"3d085a58",
  2510 => x"80568076",
  2511 => x"54547751",
  2512 => x"785281b6",
  2513 => x"fd3f8008",
  2514 => x"81a63880",
  2515 => x"c13d0858",
  2516 => x"81780c82",
  2517 => x"bcc45f8c",
  2518 => x"08802e86",
  2519 => x"38811f8c",
  2520 => x"080c7e56",
  2521 => x"75800cba",
  2522 => x"3d0d8c0c",
  2523 => x"047f80c4",
  2524 => x"05088417",
  2525 => x"0c816080",
  2526 => x"c405082b",
  2527 => x"88170c75",
  2528 => x"527f5180",
  2529 => x"c7f23f67",
  2530 => x"6080c005",
  2531 => x"0cb83d08",
  2532 => x"57768025",
  2533 => x"ff893881",
  2534 => x"7a0c76fe",
  2535 => x"0a0670ba",
  2536 => x"3d0c709f",
  2537 => x"fe0a0657",
  2538 => x"57759ffe",
  2539 => x"0a2e0981",
  2540 => x"06fefd38",
  2541 => x"80c13d08",
  2542 => x"5680ce8f",
  2543 => x"760cb93d",
  2544 => x"0883ff38",
  2545 => x"76bfffff",
  2546 => x"0682bcf8",
  2547 => x"40567583",
  2548 => x"f1388c08",
  2549 => x"802eff8a",
  2550 => x"38831f33",
  2551 => x"7f880558",
  2552 => x"56758438",
  2553 => x"831f5776",
  2554 => x"8c080c7e",
  2555 => x"56fef539",
  2556 => x"ba3dffb4",
  2557 => x"1156ffb0",
  2558 => x"05547752",
  2559 => x"78537f51",
  2560 => x"80d7933f",
  2561 => x"8008b93d",
  2562 => x"0870942a",
  2563 => x"8fff065e",
  2564 => x"59417b83",
  2565 => x"b438a73d",
  2566 => x"08a73d08",
  2567 => x"0588b211",
  2568 => x"5d56a07c",
  2569 => x"258e8138",
  2570 => x"80c07c31",
  2571 => x"88921779",
  2572 => x"722bbc3d",
  2573 => x"08722a07",
  2574 => x"b53d7156",
  2575 => x"70555d51",
  2576 => x"575781be",
  2577 => x"8f3fb23d",
  2578 => x"08b43d08",
  2579 => x"b23d5d5a",
  2580 => x"58807624",
  2581 => x"91a23877",
  2582 => x"b73d0c78",
  2583 => x"b83d0cb6",
  2584 => x"3d0890ff",
  2585 => x"0a05b73d",
  2586 => x"0cf7cd1c",
  2587 => x"5c814ebf",
  2588 => x"fc0a5680",
  2589 => x"765555b6",
  2590 => x"3d08b83d",
  2591 => x"08585276",
  2592 => x"537a5181",
  2593 => x"85d43f83",
  2594 => x"feca8fa7",
  2595 => x"56869bbd",
  2596 => x"86e17655",
  2597 => x"55b03d08",
  2598 => x"b23d0858",
  2599 => x"52765379",
  2600 => x"518186e0",
  2601 => x"3f83fe9a",
  2602 => x"94a856f8",
  2603 => x"db8391b3",
  2604 => x"765555b2",
  2605 => x"3d08b43d",
  2606 => x"08585276",
  2607 => x"53ba3dd0",
  2608 => x"05518183",
  2609 => x"f73fae3d",
  2610 => x"08b03d08",
  2611 => x"7d54ae3d",
  2612 => x"535a5881",
  2613 => x"bcfe3faa",
  2614 => x"3d4c83fe",
  2615 => x"cd889356",
  2616 => x"8584fdf3",
  2617 => x"fb765555",
  2618 => x"ac3d08ae",
  2619 => x"3d085852",
  2620 => x"76536b51",
  2621 => x"81868d3f",
  2622 => x"a83dab3d",
  2623 => x"08ad3d08",
  2624 => x"59557756",
  2625 => x"78537954",
  2626 => x"70524581",
  2627 => x"83ae3fa8",
  2628 => x"3d08aa3d",
  2629 => x"08715370",
  2630 => x"545f5d81",
  2631 => x"beb13f80",
  2632 => x"08438056",
  2633 => x"80765454",
  2634 => x"7c517d52",
  2635 => x"81b8d13f",
  2636 => x"800b8008",
  2637 => x"248cc338",
  2638 => x"810ba23d",
  2639 => x"0c629626",
  2640 => x"ae386210",
  2641 => x"101082be",
  2642 => x"ac058411",
  2643 => x"08710855",
  2644 => x"55b93d08",
  2645 => x"bb3d0859",
  2646 => x"52567652",
  2647 => x"81b8a13f",
  2648 => x"800b8008",
  2649 => x"24637131",
  2650 => x"4456800b",
  2651 => x"a23d0ca7",
  2652 => x"3d087c31",
  2653 => x"ff055a80",
  2654 => x"7a454b6a",
  2655 => x"7a248bd1",
  2656 => x"38806324",
  2657 => x"9aad3880",
  2658 => x"0ba63d0c",
  2659 => x"624f6363",
  2660 => x"05448962",
  2661 => x"27833880",
  2662 => x"42815885",
  2663 => x"62258738",
  2664 => x"61fc0542",
  2665 => x"8058810b",
  2666 => x"a13d0cff",
  2667 => x"70a53d0c",
  2668 => x"46618526",
  2669 => x"829c3861",
  2670 => x"101082bd",
  2671 => x"84055675",
  2672 => x"080482bc",
  2673 => x"cc5ffc8a",
  2674 => x"39b83d08",
  2675 => x"ba3d0858",
  2676 => x"b73d0c76",
  2677 => x"b83d0cb6",
  2678 => x"3d08fc0a",
  2679 => x"069ffc0a",
  2680 => x"07b73d0c",
  2681 => x"f8811c5c",
  2682 => x"804eb23d",
  2683 => x"b13d5c5a",
  2684 => x"bffc0a56",
  2685 => x"80765555",
  2686 => x"b63d08b8",
  2687 => x"3d085852",
  2688 => x"76537a51",
  2689 => x"8182d33f",
  2690 => x"83feca8f",
  2691 => x"a756869b",
  2692 => x"bd86e176",
  2693 => x"5555b03d",
  2694 => x"08b23d08",
  2695 => x"58527653",
  2696 => x"79518183",
  2697 => x"df3f83fe",
  2698 => x"9a94a856",
  2699 => x"f8db8391",
  2700 => x"b3765555",
  2701 => x"b23d08b4",
  2702 => x"3d085852",
  2703 => x"7653ba3d",
  2704 => x"d0055181",
  2705 => x"80f63fae",
  2706 => x"3d08b03d",
  2707 => x"087d54ae",
  2708 => x"3d535a58",
  2709 => x"81b9fd3f",
  2710 => x"aa3d4c83",
  2711 => x"fecd8893",
  2712 => x"568584fd",
  2713 => x"f3fb7655",
  2714 => x"55ac3d08",
  2715 => x"ae3d0858",
  2716 => x"5276536b",
  2717 => x"5181838c",
  2718 => x"3fa83dab",
  2719 => x"3d08ad3d",
  2720 => x"08595577",
  2721 => x"56785379",
  2722 => x"54705245",
  2723 => x"8180ad3f",
  2724 => x"a83d08aa",
  2725 => x"3d087153",
  2726 => x"70545f5d",
  2727 => x"81bbb03f",
  2728 => x"80084380",
  2729 => x"56807654",
  2730 => x"547c517d",
  2731 => x"5281b5d0",
  2732 => x"3f800880",
  2733 => x"25fd8138",
  2734 => x"89c03980",
  2735 => x"0ba13d0c",
  2736 => x"68630581",
  2737 => x"1170485d",
  2738 => x"a43d0c7b",
  2739 => x"80248338",
  2740 => x"815c845a",
  2741 => x"806080c4",
  2742 => x"050c987c",
  2743 => x"26973880",
  2744 => x"5781177a",
  2745 => x"10941158",
  2746 => x"5b577b76",
  2747 => x"27f33876",
  2748 => x"6080c405",
  2749 => x"0c7f80c4",
  2750 => x"0508527f",
  2751 => x"51bfef3f",
  2752 => x"80086080",
  2753 => x"c0050c80",
  2754 => x"0880088e",
  2755 => x"68275840",
  2756 => x"4d77802e",
  2757 => x"86903875",
  2758 => x"802e868a",
  2759 => x"38b83d08",
  2760 => x"ba3d0871",
  2761 => x"b93d0c70",
  2762 => x"ba3d0c64",
  2763 => x"a53d0c67",
  2764 => x"a73d0c5a",
  2765 => x"58825c80",
  2766 => x"63258ad7",
  2767 => x"3862832b",
  2768 => x"80f80682",
  2769 => x"beac1108",
  2770 => x"82beb012",
  2771 => x"0865842c",
  2772 => x"70842a70",
  2773 => x"81065154",
  2774 => x"5d405e56",
  2775 => x"7588e438",
  2776 => x"79802e9f",
  2777 => x"3882be84",
  2778 => x"58798106",
  2779 => x"567587e9",
  2780 => x"3879812c",
  2781 => x"8819595a",
  2782 => x"79ef38b8",
  2783 => x"3d08ba3d",
  2784 => x"085a587c",
  2785 => x"547d5577",
  2786 => x"52785364",
  2787 => x"51819e83",
  2788 => x"3fa83d08",
  2789 => x"aa3d0871",
  2790 => x"bb3d0c70",
  2791 => x"bc3d0c5a",
  2792 => x"58a13d08",
  2793 => x"802e80d9",
  2794 => x"38805a9f",
  2795 => x"fc0a5680",
  2796 => x"76545477",
  2797 => x"51785281",
  2798 => x"b3c63f79",
  2799 => x"8008248b",
  2800 => x"f3388066",
  2801 => x"25bb3879",
  2802 => x"802eb638",
  2803 => x"800ba43d",
  2804 => x"082584ba",
  2805 => x"38a33d08",
  2806 => x"63ff0544",
  2807 => x"4680c882",
  2808 => x"0a568076",
  2809 => x"55557752",
  2810 => x"78536451",
  2811 => x"8180953f",
  2812 => x"a83d08aa",
  2813 => x"3d085ab9",
  2814 => x"3d0c78ba",
  2815 => x"3d0c811c",
  2816 => x"5c7b5264",
  2817 => x"5181b6cc",
  2818 => x"3fb83d08",
  2819 => x"ba3d0858",
  2820 => x"547655a8",
  2821 => x"3d08aa3d",
  2822 => x"08585276",
  2823 => x"536b5180",
  2824 => x"ffe23f80",
  2825 => x"f0820a56",
  2826 => x"80765555",
  2827 => x"aa3d08ac",
  2828 => x"3d085852",
  2829 => x"7653ac3d",
  2830 => x"5180fd80",
  2831 => x"3fac3d08",
  2832 => x"ae3d0858",
  2833 => x"b53d0c76",
  2834 => x"b63d0cb4",
  2835 => x"3d0886bf",
  2836 => x"0a05b53d",
  2837 => x"0c65802e",
  2838 => x"96bd386f",
  2839 => x"802e94f2",
  2840 => x"38651010",
  2841 => x"1082bea4",
  2842 => x"05841108",
  2843 => x"71085656",
  2844 => x"568ffc0a",
  2845 => x"56807653",
  2846 => x"53645181",
  2847 => x"9c953fb4",
  2848 => x"3d08b63d",
  2849 => x"08585476",
  2850 => x"55a83d08",
  2851 => x"aa3d0858",
  2852 => x"5276536b",
  2853 => x"5180fdc2",
  2854 => x"3faa3d08",
  2855 => x"ac3d0858",
  2856 => x"b53d0c76",
  2857 => x"b63d0c80",
  2858 => x"0bb93d08",
  2859 => x"bb3d085b",
  2860 => x"595c80c8",
  2861 => x"820a5d80",
  2862 => x"5e775178",
  2863 => x"5281b78f",
  2864 => x"3f800880",
  2865 => x"08536552",
  2866 => x"5a81b588",
  2867 => x"3fa83d08",
  2868 => x"aa3d0858",
  2869 => x"547655b8",
  2870 => x"3d08ba3d",
  2871 => x"08585276",
  2872 => x"536b5180",
  2873 => x"fcf43faa",
  2874 => x"3d08ac3d",
  2875 => x"085ab93d",
  2876 => x"0c78ba3d",
  2877 => x"0cb01a56",
  2878 => x"757f7081",
  2879 => x"054134b8",
  2880 => x"3d08ba3d",
  2881 => x"08b63d08",
  2882 => x"b83d085a",
  2883 => x"55785671",
  2884 => x"5370545a",
  2885 => x"5881b0e8",
  2886 => x"3f800b80",
  2887 => x"082486cc",
  2888 => x"38775478",
  2889 => x"559ffc0a",
  2890 => x"56807653",
  2891 => x"53645180",
  2892 => x"fca83fb4",
  2893 => x"3d08b63d",
  2894 => x"08715570",
  2895 => x"56aa3d08",
  2896 => x"ac3d085a",
  2897 => x"5378545a",
  2898 => x"5881b0b4",
  2899 => x"3f800b80",
  2900 => x"082485ed",
  2901 => x"38811c5c",
  2902 => x"7b662581",
  2903 => x"b1387c54",
  2904 => x"7d557752",
  2905 => x"78536b51",
  2906 => x"80fd993f",
  2907 => x"aa3d08ac",
  2908 => x"3d0858b5",
  2909 => x"3d0c76b6",
  2910 => x"3d0c7c54",
  2911 => x"7d55b83d",
  2912 => x"08ba3d08",
  2913 => x"58527653",
  2914 => x"645180fc",
  2915 => x"f73fa83d",
  2916 => x"08aa3d08",
  2917 => x"71bb3d0c",
  2918 => x"70bc3d0c",
  2919 => x"5a58fe99",
  2920 => x"398ffc0a",
  2921 => x"58807855",
  2922 => x"7056b53d",
  2923 => x"08b73d08",
  2924 => x"59537754",
  2925 => x"65525980",
  2926 => x"fa823fa8",
  2927 => x"3d08aa3d",
  2928 => x"08585376",
  2929 => x"54b83d08",
  2930 => x"ba3d0858",
  2931 => x"51765281",
  2932 => x"adc43f80",
  2933 => x"08802484",
  2934 => x"e838b43d",
  2935 => x"08b63d08",
  2936 => x"58547655",
  2937 => x"77527853",
  2938 => x"6b5180fa",
  2939 => x"ed3faa3d",
  2940 => x"08ac3d08",
  2941 => x"58537654",
  2942 => x"b83d08ba",
  2943 => x"3d085851",
  2944 => x"765281ae",
  2945 => x"fb3f800b",
  2946 => x"80082492",
  2947 => x"f9386cb7",
  2948 => x"3d08b93d",
  2949 => x"085bba3d",
  2950 => x"0c79bb3d",
  2951 => x"0ca33d08",
  2952 => x"a63d0848",
  2953 => x"445f800b",
  2954 => x"a73d0857",
  2955 => x"58777624",
  2956 => x"83388158",
  2957 => x"80780657",
  2958 => x"628e2487",
  2959 => x"e5388170",
  2960 => x"79065859",
  2961 => x"76802e87",
  2962 => x"d9386210",
  2963 => x"101082be",
  2964 => x"ac057008",
  2965 => x"84120880",
  2966 => x"6c245340",
  2967 => x"5e568066",
  2968 => x"2585c838",
  2969 => x"810bb93d",
  2970 => x"08bb3d08",
  2971 => x"5b595c7c",
  2972 => x"547d5577",
  2973 => x"52785364",
  2974 => x"51819897",
  2975 => x"3fa83d08",
  2976 => x"aa3d0858",
  2977 => x"51765281",
  2978 => x"b3c53f80",
  2979 => x"08800853",
  2980 => x"65525a81",
  2981 => x"b1be3f7c",
  2982 => x"547d55a8",
  2983 => x"3d08aa3d",
  2984 => x"08585276",
  2985 => x"536b5180",
  2986 => x"fada3faa",
  2987 => x"3d08ac3d",
  2988 => x"08585476",
  2989 => x"55b83d08",
  2990 => x"ba3d0858",
  2991 => x"527653ac",
  2992 => x"3d5180f9",
  2993 => x"953fac3d",
  2994 => x"08ae3d08",
  2995 => x"5ab93d0c",
  2996 => x"78ba3d0c",
  2997 => x"b01a5675",
  2998 => x"7f708105",
  2999 => x"41347b66",
  3000 => x"2e828f38",
  3001 => x"80c8820a",
  3002 => x"56807655",
  3003 => x"55b83d08",
  3004 => x"ba3d0858",
  3005 => x"52765364",
  3006 => x"5180fa88",
  3007 => x"3fa83d08",
  3008 => x"aa3d0871",
  3009 => x"bb3d0c70",
  3010 => x"bc3d0c5a",
  3011 => x"58805680",
  3012 => x"76545477",
  3013 => x"51785281",
  3014 => x"a7a83f80",
  3015 => x"08802e82",
  3016 => x"cb38811c",
  3017 => x"5cfec839",
  3018 => x"a07c31ba",
  3019 => x"3d08712b",
  3020 => x"b43d7155",
  3021 => x"70545c51",
  3022 => x"5681b098",
  3023 => x"3fb23d08",
  3024 => x"b43d08b2",
  3025 => x"3d5d5a58",
  3026 => x"758025f2",
  3027 => x"8a3883a8",
  3028 => x"3979304b",
  3029 => x"8044f4a9",
  3030 => x"39811c78",
  3031 => x"08841a08",
  3032 => x"59557756",
  3033 => x"7d537e54",
  3034 => x"65525c80",
  3035 => x"f9963fa8",
  3036 => x"3d08aa3d",
  3037 => x"085f5df7",
  3038 => x"f8396252",
  3039 => x"645181af",
  3040 => x"d33f7c53",
  3041 => x"7d54a83d",
  3042 => x"08aa3d08",
  3043 => x"58517652",
  3044 => x"81a8993f",
  3045 => x"80083070",
  3046 => x"8008079f",
  3047 => x"2a647131",
  3048 => x"455156f3",
  3049 => x"9339800b",
  3050 => x"a13d0c80",
  3051 => x"692583f7",
  3052 => x"386869a5",
  3053 => x"3d0c6947",
  3054 => x"5cf69739",
  3055 => x"925c8049",
  3056 => x"f6903979",
  3057 => x"8f0682be",
  3058 => x"a40882be",
  3059 => x"a8085955",
  3060 => x"77567853",
  3061 => x"79546552",
  3062 => x"5a8195b7",
  3063 => x"3fa83d08",
  3064 => x"aa3d0871",
  3065 => x"bb3d0c70",
  3066 => x"bc3d0c5a",
  3067 => x"58835cf6",
  3068 => x"ef39b83d",
  3069 => x"08ba3d08",
  3070 => x"71567057",
  3071 => x"58527653",
  3072 => x"645180f5",
  3073 => x"b73fa83d",
  3074 => x"08aa3d08",
  3075 => x"71bb3d0c",
  3076 => x"70bc3d0c",
  3077 => x"7e557f56",
  3078 => x"71537054",
  3079 => x"5a5881a8",
  3080 => x"f53f8008",
  3081 => x"80249a38",
  3082 => x"7c537d54",
  3083 => x"77517852",
  3084 => x"81a58f3f",
  3085 => x"8008b538",
  3086 => x"79810656",
  3087 => x"75802eac",
  3088 => x"38ff1f70",
  3089 => x"33575f75",
  3090 => x"b92e0981",
  3091 => x"0690387e",
  3092 => x"6d2e0981",
  3093 => x"06eb3862",
  3094 => x"810543b0",
  3095 => x"6d347e7f",
  3096 => x"81057133",
  3097 => x"81055840",
  3098 => x"57757734",
  3099 => x"60527f51",
  3100 => x"b6863f80",
  3101 => x"7f3480c1",
  3102 => x"3d086381",
  3103 => x"05710c56",
  3104 => x"8c08802e",
  3105 => x"85387e8c",
  3106 => x"080c6c80",
  3107 => x"0cba3d0d",
  3108 => x"8c0c0462",
  3109 => x"305b7a80",
  3110 => x"2ef68638",
  3111 => x"7a832b80",
  3112 => x"f80682be",
  3113 => x"b0110882",
  3114 => x"beac1208",
  3115 => x"56567853",
  3116 => x"79546552",
  3117 => x"5680f6cc",
  3118 => x"3fa83d08",
  3119 => x"aa3d0871",
  3120 => x"bb3d0c70",
  3121 => x"bc3d0c7c",
  3122 => x"842c5c5a",
  3123 => x"5879802e",
  3124 => x"f5cf3882",
  3125 => x"be847a81",
  3126 => x"06575b75",
  3127 => x"81db3879",
  3128 => x"812c881c",
  3129 => x"5c5a7980",
  3130 => x"2ef5b638",
  3131 => x"79810656",
  3132 => x"75802eeb",
  3133 => x"3881c239",
  3134 => x"9f820a56",
  3135 => x"80765555",
  3136 => x"77527853",
  3137 => x"7a5180f3",
  3138 => x"b33fb03d",
  3139 => x"08b23d08",
  3140 => x"5ab73d0c",
  3141 => x"78b83d0c",
  3142 => x"b63d0890",
  3143 => x"ff0a05b7",
  3144 => x"3d0cf7cd",
  3145 => x"1c5c814e",
  3146 => x"eec53975",
  3147 => x"79065675",
  3148 => x"802efab0",
  3149 => x"38807048",
  3150 => x"4a696624",
  3151 => x"81de3880",
  3152 => x"d0820a56",
  3153 => x"80765555",
  3154 => x"7c527d53",
  3155 => x"645180f5",
  3156 => x"b33fa83d",
  3157 => x"08aa3d08",
  3158 => x"58537654",
  3159 => x"b83d08ba",
  3160 => x"3d085851",
  3161 => x"765281aa",
  3162 => x"813f6980",
  3163 => x"082581ac",
  3164 => x"386c5fb1",
  3165 => x"7f708105",
  3166 => x"41346281",
  3167 => x"05436652",
  3168 => x"7f51b3f4",
  3169 => x"3f69802e",
  3170 => x"fde23867",
  3171 => x"30706907",
  3172 => x"9f2a5156",
  3173 => x"676a2e85",
  3174 => x"387580d1",
  3175 => x"3869527f",
  3176 => x"51b3d53f",
  3177 => x"fdc63981",
  3178 => x"7071a63d",
  3179 => x"0c71485d",
  3180 => x"49f29f39",
  3181 => x"815af48a",
  3182 => x"39811c7b",
  3183 => x"08841d08",
  3184 => x"59557756",
  3185 => x"78537954",
  3186 => x"65525c80",
  3187 => x"f4b63fa8",
  3188 => x"3d08aa3d",
  3189 => x"0871bb3d",
  3190 => x"0c70bc3d",
  3191 => x"0c7b812c",
  3192 => x"881e5e5c",
  3193 => x"5a5879fe",
  3194 => x"8338f3b5",
  3195 => x"3967527f",
  3196 => x"51b3853f",
  3197 => x"69527f51",
  3198 => x"b2fe3ffc",
  3199 => x"ef397781",
  3200 => x"0a325378",
  3201 => x"5479517a",
  3202 => x"5281a6f4",
  3203 => x"3f800880",
  3204 => x"25f7fb38",
  3205 => x"79b93d0c",
  3206 => x"7aba3d0c",
  3207 => x"680943fe",
  3208 => x"dd396aa6",
  3209 => x"3d087879",
  3210 => x"4b4c5959",
  3211 => x"6f802e80",
  3212 => x"c3388162",
  3213 => x"258bb938",
  3214 => x"65ff05a6",
  3215 => x"3d087131",
  3216 => x"595aa53d",
  3217 => x"087a2594",
  3218 => x"3879a63d",
  3219 => x"08316f11",
  3220 => x"a13d0ca6",
  3221 => x"3d0805a6",
  3222 => x"3d0c7658",
  3223 => x"655c8066",
  3224 => x"2483be38",
  3225 => x"6a1c641d",
  3226 => x"454b8152",
  3227 => x"7f51b6fc",
  3228 => x"3f80084a",
  3229 => x"78802456",
  3230 => x"8064259b",
  3231 => x"3875802e",
  3232 => x"9638635c",
  3233 => x"78642583",
  3234 => x"38785c6a",
  3235 => x"7c31797d",
  3236 => x"31657e31",
  3237 => x"465a4b80",
  3238 => x"0ba63d08",
  3239 => x"25b8386f",
  3240 => x"802e889d",
  3241 => x"38807825",
  3242 => x"a3387753",
  3243 => x"69527f51",
  3244 => x"b99c3f80",
  3245 => x"08615480",
  3246 => x"08536052",
  3247 => x"4ab6c83f",
  3248 => x"80086153",
  3249 => x"605256b1",
  3250 => x"af3f7541",
  3251 => x"a53d0878",
  3252 => x"315a7982",
  3253 => x"bd388152",
  3254 => x"7f51b690",
  3255 => x"3f800847",
  3256 => x"806f258e",
  3257 => x"386e5380",
  3258 => x"08527f51",
  3259 => x"b8e03f80",
  3260 => x"08478058",
  3261 => x"81622581",
  3262 => x"d6386381",
  3263 => x"059f065c",
  3264 => x"6e81b238",
  3265 => x"7b802e85",
  3266 => x"38a07c31",
  3267 => x"5c847c25",
  3268 => x"86c438fc",
  3269 => x"1c6b1171",
  3270 => x"1b5b4c64",
  3271 => x"0544806b",
  3272 => x"258d386a",
  3273 => x"5360527f",
  3274 => x"51b9e33f",
  3275 => x"80084180",
  3276 => x"64258d38",
  3277 => x"63536652",
  3278 => x"7f51b9d2",
  3279 => x"3f800847",
  3280 => x"a13d0880",
  3281 => x"c5388066",
  3282 => x"25568262",
  3283 => x"2581ff38",
  3284 => x"75802e81",
  3285 => x"f9388066",
  3286 => x"24fdc138",
  3287 => x"80548553",
  3288 => x"66527f51",
  3289 => x"b0b43f80",
  3290 => x"08800853",
  3291 => x"615247ba",
  3292 => x"e13f800b",
  3293 => x"800825fd",
  3294 => x"a3386c5f",
  3295 => x"b17f7081",
  3296 => x"05413462",
  3297 => x"810543fb",
  3298 => x"f5396652",
  3299 => x"6051bac2",
  3300 => x"3f800880",
  3301 => x"25ffaf38",
  3302 => x"62ff0543",
  3303 => x"80548a53",
  3304 => x"60527f51",
  3305 => x"aff43f80",
  3306 => x"08416f81",
  3307 => x"8c38a33d",
  3308 => x"0846ff92",
  3309 => x"39669005",
  3310 => x"08101067",
  3311 => x"05901108",
  3312 => x"5256b295",
  3313 => x"3f638008",
  3314 => x"319f065c",
  3315 => x"feb639b9",
  3316 => x"3d08782e",
  3317 => x"098106fe",
  3318 => x"a138b83d",
  3319 => x"0870bfff",
  3320 => x"ff065757",
  3321 => x"75782e09",
  3322 => x"8106fe8e",
  3323 => x"38769ffe",
  3324 => x"0a065675",
  3325 => x"782efe82",
  3326 => x"386a8105",
  3327 => x"64810545",
  3328 => x"4b816481",
  3329 => x"059f065d",
  3330 => x"586e802e",
  3331 => x"fdf638ff",
  3332 => x"a4397953",
  3333 => x"60527f51",
  3334 => x"b6b43f80",
  3335 => x"0841fdb6",
  3336 => x"396a6631",
  3337 => x"59806b11",
  3338 => x"4c640544",
  3339 => x"81527f51",
  3340 => x"b3ba3f80",
  3341 => x"084afcbc",
  3342 => x"3980548a",
  3343 => x"5369527f",
  3344 => x"51aed73f",
  3345 => x"8008a43d",
  3346 => x"08474afd",
  3347 => x"f939815c",
  3348 => x"6f802e81",
  3349 => x"ef388079",
  3350 => x"258d3878",
  3351 => x"5369527f",
  3352 => x"51b7ab3f",
  3353 => x"80084a69",
  3354 => x"48778294",
  3355 => x"38815c66",
  3356 => x"526051e2",
  3357 => x"a03f8008",
  3358 => x"b0056853",
  3359 => x"615257b8",
  3360 => x"d13f8008",
  3361 => x"6a546753",
  3362 => x"60525ab9",
  3363 => x"9c3f8008",
  3364 => x"56815b80",
  3365 => x"088c0508",
  3366 => x"802e81d6",
  3367 => x"3875527f",
  3368 => x"51add53f",
  3369 => x"7a620756",
  3370 => x"758d38b9",
  3371 => x"3d088106",
  3372 => x"5675802e",
  3373 => x"81fe3880",
  3374 => x"7a24828c",
  3375 => x"38796207",
  3376 => x"56758d38",
  3377 => x"b93d0881",
  3378 => x"06567580",
  3379 => x"2e81f938",
  3380 => x"7a802486",
  3381 => x"bc38767f",
  3382 => x"70810541",
  3383 => x"347b662e",
  3384 => x"83883880",
  3385 => x"548a5360",
  3386 => x"527f51ad",
  3387 => x"ad3f8008",
  3388 => x"41676a2e",
  3389 => x"82c93880",
  3390 => x"548a5367",
  3391 => x"527f51ad",
  3392 => x"993f8008",
  3393 => x"4880548a",
  3394 => x"5369527f",
  3395 => x"51ad8b3f",
  3396 => x"8008811d",
  3397 => x"5d4a6652",
  3398 => x"6051e0f9",
  3399 => x"3f8008b0",
  3400 => x"05685361",
  3401 => x"5257b7aa",
  3402 => x"3f80086a",
  3403 => x"54675360",
  3404 => x"525ab7f5",
  3405 => x"3f800856",
  3406 => x"815b8008",
  3407 => x"8c0508fe",
  3408 => x"dc38af39",
  3409 => x"66527e7f",
  3410 => x"81056253",
  3411 => x"4056e0c5",
  3412 => x"3f8008b0",
  3413 => x"05577676",
  3414 => x"347b6625",
  3415 => x"828c3880",
  3416 => x"548a5360",
  3417 => x"527f51ac",
  3418 => x"b13f8008",
  3419 => x"811d5d41",
  3420 => x"d3398008",
  3421 => x"526051b6",
  3422 => x"d93f8008",
  3423 => x"5bfe9e39",
  3424 => x"69840508",
  3425 => x"527f51aa",
  3426 => x"e53f8008",
  3427 => x"68900508",
  3428 => x"10108805",
  3429 => x"54688c05",
  3430 => x"5380088c",
  3431 => x"05524aff",
  3432 => x"a6ed3f81",
  3433 => x"5369527f",
  3434 => x"51b4e33f",
  3435 => x"80084a81",
  3436 => x"5cfdbc39",
  3437 => x"76b92ebb",
  3438 => x"38798024",
  3439 => x"1757767f",
  3440 => x"70810541",
  3441 => x"34f7b739",
  3442 => x"807b25f2",
  3443 => x"38815360",
  3444 => x"527f51b4",
  3445 => x"b93f8008",
  3446 => x"67538008",
  3447 => x"5241b5f2",
  3448 => x"3f800b80",
  3449 => x"0825ba38",
  3450 => x"81175776",
  3451 => x"ba2e0981",
  3452 => x"06cc38b9",
  3453 => x"7f708105",
  3454 => x"4134ff1f",
  3455 => x"7033575f",
  3456 => x"75b92e09",
  3457 => x"8106819a",
  3458 => x"387e6d2e",
  3459 => x"098106ea",
  3460 => x"38628105",
  3461 => x"6d4043b1",
  3462 => x"7f708105",
  3463 => x"4134f6de",
  3464 => x"398008ff",
  3465 => x"99387681",
  3466 => x"06567580",
  3467 => x"2eff8f38",
  3468 => x"81175776",
  3469 => x"ba2e0981",
  3470 => x"06ff8338",
  3471 => x"ffb53980",
  3472 => x"548a5369",
  3473 => x"527f51aa",
  3474 => x"d13f8008",
  3475 => x"8008811e",
  3476 => x"5e494afd",
  3477 => x"c1397b83",
  3478 => x"24f9c338",
  3479 => x"9c1c6b11",
  3480 => x"711b5b4c",
  3481 => x"640544f9",
  3482 => x"b5398153",
  3483 => x"60527f51",
  3484 => x"b39c3f80",
  3485 => x"08675380",
  3486 => x"085241b4",
  3487 => x"d53f8008",
  3488 => x"8024fef6",
  3489 => x"38800889",
  3490 => x"38768106",
  3491 => x"5675feea",
  3492 => x"38ff1f70",
  3493 => x"33575f75",
  3494 => x"b02ef638",
  3495 => x"811f5ff5",
  3496 => x"dd397e7f",
  3497 => x"81057133",
  3498 => x"81055840",
  3499 => x"57757734",
  3500 => x"f5cc396a",
  3501 => x"63316330",
  3502 => x"a73d0c4b",
  3503 => x"804fe5d2",
  3504 => x"39a53d08",
  3505 => x"5360527f",
  3506 => x"51b1833f",
  3507 => x"800841f8",
  3508 => x"85396510",
  3509 => x"101082be",
  3510 => x"a4058411",
  3511 => x"08710856",
  3512 => x"56b53d08",
  3513 => x"b73d0859",
  3514 => x"53567653",
  3515 => x"645180ea",
  3516 => x"933fa83d",
  3517 => x"08aa3d08",
  3518 => x"58b53d0c",
  3519 => x"76b63d0c",
  3520 => x"810bb93d",
  3521 => x"08bb3d08",
  3522 => x"5b595c77",
  3523 => x"51785281",
  3524 => x"a2bd3f80",
  3525 => x"08800853",
  3526 => x"65525a81",
  3527 => x"a0b63fa8",
  3528 => x"3d08aa3d",
  3529 => x"08585476",
  3530 => x"55b83d08",
  3531 => x"ba3d0858",
  3532 => x"5276536b",
  3533 => x"5180e8a2",
  3534 => x"3faa3d08",
  3535 => x"ac3d085a",
  3536 => x"b93d0c78",
  3537 => x"ba3d0cb0",
  3538 => x"1a56757f",
  3539 => x"70810541",
  3540 => x"347b662e",
  3541 => x"eccb3881",
  3542 => x"1c5c80c8",
  3543 => x"820a5680",
  3544 => x"765555b8",
  3545 => x"3d08ba3d",
  3546 => x"08585276",
  3547 => x"53645180",
  3548 => x"e9923fa8",
  3549 => x"3d08aa3d",
  3550 => x"0871bb3d",
  3551 => x"0c70bc3d",
  3552 => x"0c5a58ff",
  3553 => x"8639ff1f",
  3554 => x"7033575f",
  3555 => x"75b02ef6",
  3556 => x"38811f5f",
  3557 => x"f1d63965",
  3558 => x"66484a80",
  3559 => x"d0820a56",
  3560 => x"80765555",
  3561 => x"b83d08ba",
  3562 => x"3d085852",
  3563 => x"76536451",
  3564 => x"80e7a73f",
  3565 => x"a83d08aa",
  3566 => x"3d08b63d",
  3567 => x"08b83d08",
  3568 => x"71577058",
  3569 => x"73557256",
  3570 => x"5c5a5c5a",
  3571 => x"8199c73f",
  3572 => x"800b8008",
  3573 => x"25f4a738",
  3574 => x"79b93d0c",
  3575 => x"7aba3d0c",
  3576 => x"6c5fb17f",
  3577 => x"70810541",
  3578 => x"34628105",
  3579 => x"43f38f39",
  3580 => x"88b3165c",
  3581 => x"6df4ed38",
  3582 => x"b60ba83d",
  3583 => x"08316b11",
  3584 => x"4c640544",
  3585 => x"81527f51",
  3586 => x"abe23f80",
  3587 => x"084af4e4",
  3588 => x"3976b92e",
  3589 => x"fbdd3881",
  3590 => x"1756757f",
  3591 => x"70810541",
  3592 => x"34f2db39",
  3593 => x"f83d0d7a",
  3594 => x"5877802e",
  3595 => x"81993882",
  3596 => x"c0c00854",
  3597 => x"b8140880",
  3598 => x"2e80ed38",
  3599 => x"8c182270",
  3600 => x"902b7090",
  3601 => x"2c70832a",
  3602 => x"81328106",
  3603 => x"5c515754",
  3604 => x"7880cd38",
  3605 => x"90180857",
  3606 => x"76802e80",
  3607 => x"c3387708",
  3608 => x"77317779",
  3609 => x"0c768306",
  3610 => x"7a585555",
  3611 => x"73853894",
  3612 => x"18085675",
  3613 => x"88190c80",
  3614 => x"7525a538",
  3615 => x"74537652",
  3616 => x"9c180851",
  3617 => x"a4180854",
  3618 => x"732d800b",
  3619 => x"80082580",
  3620 => x"ca388008",
  3621 => x"17758008",
  3622 => x"31565774",
  3623 => x"8024dd38",
  3624 => x"800b800c",
  3625 => x"8a3d0d04",
  3626 => x"735181db",
  3627 => x"3f8c1822",
  3628 => x"70902b70",
  3629 => x"902c7083",
  3630 => x"2a813281",
  3631 => x"065c5157",
  3632 => x"5478dd38",
  3633 => x"ff8e3980",
  3634 => x"f0a45282",
  3635 => x"c0c00851",
  3636 => x"8fdc3f80",
  3637 => x"08800c8a",
  3638 => x"3d0d048c",
  3639 => x"182280c0",
  3640 => x"0754738c",
  3641 => x"1923ff0b",
  3642 => x"800c8a3d",
  3643 => x"0d04803d",
  3644 => x"0d725180",
  3645 => x"710c800b",
  3646 => x"84120c80",
  3647 => x"0b88120c",
  3648 => x"028e0522",
  3649 => x"8c122302",
  3650 => x"9205228e",
  3651 => x"1223800b",
  3652 => x"90120c80",
  3653 => x"0b94120c",
  3654 => x"800b9812",
  3655 => x"0c709c12",
  3656 => x"0c81b7bf",
  3657 => x"0ba0120c",
  3658 => x"81b88b0b",
  3659 => x"a4120c81",
  3660 => x"b9870ba8",
  3661 => x"120c81b9",
  3662 => x"d80bac12",
  3663 => x"0c823d0d",
  3664 => x"04fa3d0d",
  3665 => x"797080dc",
  3666 => x"298c1154",
  3667 => x"7a535657",
  3668 => x"93b33f80",
  3669 => x"08800855",
  3670 => x"56800880",
  3671 => x"2ea23880",
  3672 => x"088c0554",
  3673 => x"800b8008",
  3674 => x"0c768008",
  3675 => x"84050c73",
  3676 => x"80088805",
  3677 => x"0c745380",
  3678 => x"527351a1",
  3679 => x"e03f7554",
  3680 => x"73800c88",
  3681 => x"3d0d04fc",
  3682 => x"3d0d7680",
  3683 => x"f59b0bbc",
  3684 => x"120c5581",
  3685 => x"0bb8160c",
  3686 => x"800b84dc",
  3687 => x"160c830b",
  3688 => x"84e0160c",
  3689 => x"84e81584",
  3690 => x"e4160c74",
  3691 => x"54805384",
  3692 => x"52841508",
  3693 => x"51feb73f",
  3694 => x"74548153",
  3695 => x"89528815",
  3696 => x"0851feaa",
  3697 => x"3f745482",
  3698 => x"538a528c",
  3699 => x"150851fe",
  3700 => x"9d3f863d",
  3701 => x"0d04f93d",
  3702 => x"0d7982c0",
  3703 => x"c0085457",
  3704 => x"b8130880",
  3705 => x"2e80c838",
  3706 => x"84dc1356",
  3707 => x"88160884",
  3708 => x"1708ff05",
  3709 => x"55558074",
  3710 => x"249f388c",
  3711 => x"15227090",
  3712 => x"2b70902c",
  3713 => x"51545872",
  3714 => x"802e80ca",
  3715 => x"3880dc15",
  3716 => x"ff155555",
  3717 => x"738025e3",
  3718 => x"38750853",
  3719 => x"72802e9f",
  3720 => x"38725688",
  3721 => x"16088417",
  3722 => x"08ff0555",
  3723 => x"55c83972",
  3724 => x"51fed43f",
  3725 => x"82c0c008",
  3726 => x"84dc0556",
  3727 => x"ffae3984",
  3728 => x"527651fd",
  3729 => x"fc3f8008",
  3730 => x"760c8008",
  3731 => x"802e80c0",
  3732 => x"38800856",
  3733 => x"ce39810b",
  3734 => x"8c162372",
  3735 => x"750c7288",
  3736 => x"160c7284",
  3737 => x"160c7290",
  3738 => x"160c7294",
  3739 => x"160c7298",
  3740 => x"160cff0b",
  3741 => x"8e162372",
  3742 => x"b0160c72",
  3743 => x"b4160c72",
  3744 => x"80c4160c",
  3745 => x"7280c816",
  3746 => x"0c74800c",
  3747 => x"893d0d04",
  3748 => x"8c770c80",
  3749 => x"0b800c89",
  3750 => x"3d0d04ff",
  3751 => x"3d0d80f0",
  3752 => x"a4527351",
  3753 => x"8c883f83",
  3754 => x"3d0d0480",
  3755 => x"3d0d82c0",
  3756 => x"c00851e7",
  3757 => x"3f823d0d",
  3758 => x"04fb3d0d",
  3759 => x"77705256",
  3760 => x"a0aa3f82",
  3761 => x"c89c0b88",
  3762 => x"05088411",
  3763 => x"08fc0670",
  3764 => x"7b319fef",
  3765 => x"05e08006",
  3766 => x"e0800556",
  3767 => x"5653a080",
  3768 => x"74249538",
  3769 => x"80527551",
  3770 => x"80c0c93f",
  3771 => x"82c8a408",
  3772 => x"15537280",
  3773 => x"082e8f38",
  3774 => x"75519ff1",
  3775 => x"3f805372",
  3776 => x"800c873d",
  3777 => x"0d047330",
  3778 => x"52755180",
  3779 => x"c0a63f80",
  3780 => x"08ff2ea8",
  3781 => x"3882c89c",
  3782 => x"0b880508",
  3783 => x"75753181",
  3784 => x"0784120c",
  3785 => x"5382c7e0",
  3786 => x"08743182",
  3787 => x"c7e00c75",
  3788 => x"519fba3f",
  3789 => x"810b800c",
  3790 => x"873d0d04",
  3791 => x"80527551",
  3792 => x"bff23f82",
  3793 => x"c89c0b88",
  3794 => x"05088008",
  3795 => x"71315653",
  3796 => x"8f7525ff",
  3797 => x"a3388008",
  3798 => x"82c89008",
  3799 => x"3182c7e0",
  3800 => x"0c748107",
  3801 => x"84140c75",
  3802 => x"519f823f",
  3803 => x"8053ff8f",
  3804 => x"39f63d0d",
  3805 => x"7c7e545b",
  3806 => x"72802e82",
  3807 => x"83387a51",
  3808 => x"9eea3ff8",
  3809 => x"13841108",
  3810 => x"70fe0670",
  3811 => x"13841108",
  3812 => x"fc065d58",
  3813 => x"59545882",
  3814 => x"c8a40875",
  3815 => x"2e82de38",
  3816 => x"7884160c",
  3817 => x"80738106",
  3818 => x"545a727a",
  3819 => x"2e81d538",
  3820 => x"78158411",
  3821 => x"08810651",
  3822 => x"5372a038",
  3823 => x"78175779",
  3824 => x"81e63888",
  3825 => x"15085372",
  3826 => x"82c8a42e",
  3827 => x"82f9388c",
  3828 => x"1508708c",
  3829 => x"150c7388",
  3830 => x"120c5676",
  3831 => x"81078419",
  3832 => x"0c761877",
  3833 => x"710c5379",
  3834 => x"81913883",
  3835 => x"ff772781",
  3836 => x"c8387689",
  3837 => x"2a77832a",
  3838 => x"56537280",
  3839 => x"2ebf3876",
  3840 => x"862ab805",
  3841 => x"55847327",
  3842 => x"b43880db",
  3843 => x"13559473",
  3844 => x"27ab3876",
  3845 => x"8c2a80ee",
  3846 => x"055580d4",
  3847 => x"73279e38",
  3848 => x"768f2a80",
  3849 => x"f7055582",
  3850 => x"d4732791",
  3851 => x"3876922a",
  3852 => x"80fc0555",
  3853 => x"8ad47327",
  3854 => x"843880fe",
  3855 => x"55741010",
  3856 => x"1082c89c",
  3857 => x"05881108",
  3858 => x"55567376",
  3859 => x"2e82b338",
  3860 => x"841408fc",
  3861 => x"06537673",
  3862 => x"278d3888",
  3863 => x"14085473",
  3864 => x"762e0981",
  3865 => x"06ea388c",
  3866 => x"1408708c",
  3867 => x"1a0c7488",
  3868 => x"1a0c7888",
  3869 => x"120c5677",
  3870 => x"8c150c7a",
  3871 => x"519cee3f",
  3872 => x"8c3d0d04",
  3873 => x"77087871",
  3874 => x"31597705",
  3875 => x"88190854",
  3876 => x"577282c8",
  3877 => x"a42e80e0",
  3878 => x"388c1808",
  3879 => x"708c150c",
  3880 => x"7388120c",
  3881 => x"56fe8939",
  3882 => x"8815088c",
  3883 => x"1608708c",
  3884 => x"130c5788",
  3885 => x"170cfea3",
  3886 => x"3976832a",
  3887 => x"70545580",
  3888 => x"75248198",
  3889 => x"3872822c",
  3890 => x"81712b82",
  3891 => x"c8a00807",
  3892 => x"82c89c0b",
  3893 => x"84050c53",
  3894 => x"74101010",
  3895 => x"82c89c05",
  3896 => x"88110855",
  3897 => x"56758c19",
  3898 => x"0c738819",
  3899 => x"0c778817",
  3900 => x"0c778c15",
  3901 => x"0cff8439",
  3902 => x"815afdb4",
  3903 => x"39781773",
  3904 => x"81065457",
  3905 => x"72983877",
  3906 => x"08787131",
  3907 => x"5977058c",
  3908 => x"1908881a",
  3909 => x"08718c12",
  3910 => x"0c88120c",
  3911 => x"57577681",
  3912 => x"0784190c",
  3913 => x"7782c89c",
  3914 => x"0b88050c",
  3915 => x"82c89808",
  3916 => x"7726fec7",
  3917 => x"3882c894",
  3918 => x"08527a51",
  3919 => x"fafb3f7a",
  3920 => x"519baa3f",
  3921 => x"feba3981",
  3922 => x"788c150c",
  3923 => x"7888150c",
  3924 => x"738c1a0c",
  3925 => x"73881a0c",
  3926 => x"5afd8039",
  3927 => x"83157082",
  3928 => x"2c81712b",
  3929 => x"82c8a008",
  3930 => x"0782c89c",
  3931 => x"0b84050c",
  3932 => x"51537410",
  3933 => x"101082c8",
  3934 => x"9c058811",
  3935 => x"085556fe",
  3936 => x"e4397453",
  3937 => x"807524a7",
  3938 => x"3872822c",
  3939 => x"81712b82",
  3940 => x"c8a00807",
  3941 => x"82c89c0b",
  3942 => x"84050c53",
  3943 => x"758c190c",
  3944 => x"7388190c",
  3945 => x"7788170c",
  3946 => x"778c150c",
  3947 => x"fdcd3983",
  3948 => x"1570822c",
  3949 => x"81712b82",
  3950 => x"c8a00807",
  3951 => x"82c89c0b",
  3952 => x"84050c51",
  3953 => x"53d639f2",
  3954 => x"3d0d6062",
  3955 => x"88110870",
  3956 => x"57575f5a",
  3957 => x"74802e81",
  3958 => x"90388c1a",
  3959 => x"2270832a",
  3960 => x"81327081",
  3961 => x"06515558",
  3962 => x"73863890",
  3963 => x"1a089138",
  3964 => x"7951cdbd",
  3965 => x"3fff5480",
  3966 => x"0880ee38",
  3967 => x"8c1a2258",
  3968 => x"7d085780",
  3969 => x"7883ffff",
  3970 => x"06700a10",
  3971 => x"0a708106",
  3972 => x"51565755",
  3973 => x"73752e80",
  3974 => x"d7387490",
  3975 => x"38760884",
  3976 => x"18088819",
  3977 => x"59565974",
  3978 => x"802ef238",
  3979 => x"74548880",
  3980 => x"75278438",
  3981 => x"88805473",
  3982 => x"5378529c",
  3983 => x"1a0851a4",
  3984 => x"1a085473",
  3985 => x"2d800b80",
  3986 => x"082582e6",
  3987 => x"38800819",
  3988 => x"75800831",
  3989 => x"7f880508",
  3990 => x"80083170",
  3991 => x"6188050c",
  3992 => x"56565973",
  3993 => x"ffb43880",
  3994 => x"5473800c",
  3995 => x"903d0d04",
  3996 => x"75813270",
  3997 => x"81067641",
  3998 => x"51547380",
  3999 => x"2e81c138",
  4000 => x"74903876",
  4001 => x"08841808",
  4002 => x"88195956",
  4003 => x"5974802e",
  4004 => x"f238881a",
  4005 => x"087883ff",
  4006 => x"ff067089",
  4007 => x"2a708106",
  4008 => x"51565956",
  4009 => x"73802e82",
  4010 => x"fa387575",
  4011 => x"278d3877",
  4012 => x"872a7081",
  4013 => x"06515473",
  4014 => x"82b53874",
  4015 => x"76278338",
  4016 => x"74567553",
  4017 => x"78527908",
  4018 => x"5195cf3f",
  4019 => x"881a0876",
  4020 => x"31881b0c",
  4021 => x"7908167a",
  4022 => x"0c745675",
  4023 => x"19757731",
  4024 => x"7f880508",
  4025 => x"78317061",
  4026 => x"88050c56",
  4027 => x"56597380",
  4028 => x"2efef438",
  4029 => x"8c1a2258",
  4030 => x"ff863977",
  4031 => x"78547953",
  4032 => x"7b525695",
  4033 => x"953f881a",
  4034 => x"08783188",
  4035 => x"1b0c7908",
  4036 => x"187a0c7c",
  4037 => x"76315d7c",
  4038 => x"8e387951",
  4039 => x"f2863f80",
  4040 => x"08818f38",
  4041 => x"80085f75",
  4042 => x"19757731",
  4043 => x"7f880508",
  4044 => x"78317061",
  4045 => x"88050c56",
  4046 => x"56597380",
  4047 => x"2efea838",
  4048 => x"74818338",
  4049 => x"76088418",
  4050 => x"08881959",
  4051 => x"56597480",
  4052 => x"2ef23874",
  4053 => x"538a5278",
  4054 => x"5193a03f",
  4055 => x"80087931",
  4056 => x"81055d80",
  4057 => x"08843881",
  4058 => x"155d815f",
  4059 => x"7c58747d",
  4060 => x"27833874",
  4061 => x"58941a08",
  4062 => x"881b0811",
  4063 => x"575c807a",
  4064 => x"085c5490",
  4065 => x"1a087b27",
  4066 => x"83388154",
  4067 => x"75782584",
  4068 => x"3873ba38",
  4069 => x"7b7824fe",
  4070 => x"e2387b53",
  4071 => x"78529c1a",
  4072 => x"0851a41a",
  4073 => x"0854732d",
  4074 => x"80085680",
  4075 => x"088024fe",
  4076 => x"e2388c1a",
  4077 => x"2280c007",
  4078 => x"54738c1b",
  4079 => x"23ff5473",
  4080 => x"800c903d",
  4081 => x"0d047eff",
  4082 => x"a338ff87",
  4083 => x"39755378",
  4084 => x"527a5193",
  4085 => x"c53f7908",
  4086 => x"167a0c79",
  4087 => x"51f0c53f",
  4088 => x"8008cf38",
  4089 => x"7c76315d",
  4090 => x"7cfebc38",
  4091 => x"feac3990",
  4092 => x"1a087a08",
  4093 => x"71317611",
  4094 => x"70565a57",
  4095 => x"5282c0c0",
  4096 => x"0851aafa",
  4097 => x"3f800880",
  4098 => x"2effa738",
  4099 => x"8008901b",
  4100 => x"0c800816",
  4101 => x"7a0c7794",
  4102 => x"1b0c7488",
  4103 => x"1b0c7456",
  4104 => x"fd993979",
  4105 => x"0858901a",
  4106 => x"08782783",
  4107 => x"38815475",
  4108 => x"75278438",
  4109 => x"73b33894",
  4110 => x"1a085675",
  4111 => x"752680d3",
  4112 => x"38755378",
  4113 => x"529c1a08",
  4114 => x"51a41a08",
  4115 => x"54732d80",
  4116 => x"08568008",
  4117 => x"8024fd83",
  4118 => x"388c1a22",
  4119 => x"80c00754",
  4120 => x"738c1b23",
  4121 => x"ff54fed7",
  4122 => x"39755378",
  4123 => x"52775192",
  4124 => x"a93f7908",
  4125 => x"167a0c79",
  4126 => x"51efa93f",
  4127 => x"8008802e",
  4128 => x"fcd9388c",
  4129 => x"1a2280c0",
  4130 => x"0754738c",
  4131 => x"1b23ff54",
  4132 => x"fead3974",
  4133 => x"75547953",
  4134 => x"78525691",
  4135 => x"fd3f881a",
  4136 => x"08753188",
  4137 => x"1b0c7908",
  4138 => x"157a0cfc",
  4139 => x"ae39f93d",
  4140 => x"0d797b58",
  4141 => x"53800b82",
  4142 => x"c0c00853",
  4143 => x"5672722e",
  4144 => x"80c03884",
  4145 => x"dc135574",
  4146 => x"762eb738",
  4147 => x"88150884",
  4148 => x"1608ff05",
  4149 => x"54548073",
  4150 => x"249d388c",
  4151 => x"14227090",
  4152 => x"2b70902c",
  4153 => x"51535871",
  4154 => x"80d83880",
  4155 => x"dc14ff14",
  4156 => x"54547280",
  4157 => x"25e53874",
  4158 => x"085574d0",
  4159 => x"3882c0c0",
  4160 => x"085284dc",
  4161 => x"12557480",
  4162 => x"2eb13888",
  4163 => x"15088416",
  4164 => x"08ff0554",
  4165 => x"54807324",
  4166 => x"9c388c14",
  4167 => x"2270902b",
  4168 => x"70902c51",
  4169 => x"535871ad",
  4170 => x"3880dc14",
  4171 => x"ff145454",
  4172 => x"728025e6",
  4173 => x"38740855",
  4174 => x"74d13875",
  4175 => x"800c893d",
  4176 => x"0d047351",
  4177 => x"762d7580",
  4178 => x"080780dc",
  4179 => x"15ff1555",
  4180 => x"5556ff9e",
  4181 => x"39735176",
  4182 => x"2d758008",
  4183 => x"0780dc15",
  4184 => x"ff155555",
  4185 => x"56ca39fc",
  4186 => x"3d0d7679",
  4187 => x"55557380",
  4188 => x"2e963882",
  4189 => x"bd9c5273",
  4190 => x"51b6fa3f",
  4191 => x"80089438",
  4192 => x"77b0160c",
  4193 => x"73b4160c",
  4194 => x"82bd9c53",
  4195 => x"72800c86",
  4196 => x"3d0d0482",
  4197 => x"bcc05273",
  4198 => x"51b6da3f",
  4199 => x"80538008",
  4200 => x"732e0981",
  4201 => x"06e63877",
  4202 => x"b0160c73",
  4203 => x"b4160cd8",
  4204 => x"3982c7dc",
  4205 => x"08800c04",
  4206 => x"82bdac0b",
  4207 => x"800c04fe",
  4208 => x"3d0d7553",
  4209 => x"745282c0",
  4210 => x"c00851ff",
  4211 => x"9a3f843d",
  4212 => x"0d04803d",
  4213 => x"0d82c0c0",
  4214 => x"0851dd3f",
  4215 => x"823d0d04",
  4216 => x"ea3d0d68",
  4217 => x"8c112270",
  4218 => x"0a100a81",
  4219 => x"06575856",
  4220 => x"7480e438",
  4221 => x"8e162270",
  4222 => x"902b7090",
  4223 => x"2c515558",
  4224 => x"807424b1",
  4225 => x"38983dc4",
  4226 => x"05537352",
  4227 => x"82c0c008",
  4228 => x"51b9d23f",
  4229 => x"800b8008",
  4230 => x"24973879",
  4231 => x"83e08006",
  4232 => x"547380c0",
  4233 => x"802e8190",
  4234 => x"38738280",
  4235 => x"802e8192",
  4236 => x"388c1622",
  4237 => x"57769080",
  4238 => x"0754738c",
  4239 => x"17238880",
  4240 => x"5282c0c0",
  4241 => x"085181bd",
  4242 => x"3f80089d",
  4243 => x"388c1622",
  4244 => x"82075473",
  4245 => x"8c172380",
  4246 => x"c3167077",
  4247 => x"0c90170c",
  4248 => x"810b9417",
  4249 => x"0c983d0d",
  4250 => x"0482c0c0",
  4251 => x"0880f59b",
  4252 => x"0bbc120c",
  4253 => x"548c1622",
  4254 => x"81800754",
  4255 => x"738c1723",
  4256 => x"8008760c",
  4257 => x"80089017",
  4258 => x"0c88800b",
  4259 => x"94170c74",
  4260 => x"802ed238",
  4261 => x"8e162270",
  4262 => x"902b7090",
  4263 => x"2c535558",
  4264 => x"bfda3f80",
  4265 => x"08802eff",
  4266 => x"bc388c16",
  4267 => x"22810754",
  4268 => x"738c1723",
  4269 => x"983d0d04",
  4270 => x"810b8c17",
  4271 => x"225855fe",
  4272 => x"f439a816",
  4273 => x"0881b987",
  4274 => x"2e098106",
  4275 => x"fee3388c",
  4276 => x"16228880",
  4277 => x"0754738c",
  4278 => x"17238880",
  4279 => x"0b80cc17",
  4280 => x"0cfedb39",
  4281 => x"ff3d0d73",
  4282 => x"5282c0c0",
  4283 => x"0851963f",
  4284 => x"833d0d04",
  4285 => x"ff3d0d73",
  4286 => x"5282c0c0",
  4287 => x"0851f0f1",
  4288 => x"3f833d0d",
  4289 => x"04f33d0d",
  4290 => x"7f618b11",
  4291 => x"70f8065c",
  4292 => x"55555e72",
  4293 => x"96268338",
  4294 => x"90598079",
  4295 => x"24747a26",
  4296 => x"07538054",
  4297 => x"72742e09",
  4298 => x"810680cb",
  4299 => x"387d518f",
  4300 => x"bb3f7883",
  4301 => x"f72680c6",
  4302 => x"3878832a",
  4303 => x"70101010",
  4304 => x"82c89c05",
  4305 => x"8c110859",
  4306 => x"595a7678",
  4307 => x"2e83b038",
  4308 => x"841708fc",
  4309 => x"06568c17",
  4310 => x"08881808",
  4311 => x"718c120c",
  4312 => x"88120c58",
  4313 => x"75178411",
  4314 => x"08810784",
  4315 => x"120c537d",
  4316 => x"518efa3f",
  4317 => x"88175473",
  4318 => x"800c8f3d",
  4319 => x"0d047889",
  4320 => x"2a79832a",
  4321 => x"5b537280",
  4322 => x"2ebf3878",
  4323 => x"862ab805",
  4324 => x"5a847327",
  4325 => x"b43880db",
  4326 => x"135a9473",
  4327 => x"27ab3878",
  4328 => x"8c2a80ee",
  4329 => x"055a80d4",
  4330 => x"73279e38",
  4331 => x"788f2a80",
  4332 => x"f7055a82",
  4333 => x"d4732791",
  4334 => x"3878922a",
  4335 => x"80fc055a",
  4336 => x"8ad47327",
  4337 => x"843880fe",
  4338 => x"5a791010",
  4339 => x"1082c89c",
  4340 => x"058c1108",
  4341 => x"58557675",
  4342 => x"2ea33884",
  4343 => x"1708fc06",
  4344 => x"707a3155",
  4345 => x"56738f24",
  4346 => x"88d53873",
  4347 => x"8025fee6",
  4348 => x"388c1708",
  4349 => x"5776752e",
  4350 => x"098106df",
  4351 => x"38811a5a",
  4352 => x"82c8ac08",
  4353 => x"577682c8",
  4354 => x"a42e82c0",
  4355 => x"38841708",
  4356 => x"fc06707a",
  4357 => x"31555673",
  4358 => x"8f2481f9",
  4359 => x"3882c8a4",
  4360 => x"0b82c8b0",
  4361 => x"0c82c8a4",
  4362 => x"0b82c8ac",
  4363 => x"0c738025",
  4364 => x"feb23883",
  4365 => x"ff762783",
  4366 => x"df387589",
  4367 => x"2a76832a",
  4368 => x"55537280",
  4369 => x"2ebf3875",
  4370 => x"862ab805",
  4371 => x"54847327",
  4372 => x"b43880db",
  4373 => x"13549473",
  4374 => x"27ab3875",
  4375 => x"8c2a80ee",
  4376 => x"055480d4",
  4377 => x"73279e38",
  4378 => x"758f2a80",
  4379 => x"f7055482",
  4380 => x"d4732791",
  4381 => x"3875922a",
  4382 => x"80fc0554",
  4383 => x"8ad47327",
  4384 => x"843880fe",
  4385 => x"54731010",
  4386 => x"1082c89c",
  4387 => x"05881108",
  4388 => x"56587478",
  4389 => x"2e86cf38",
  4390 => x"841508fc",
  4391 => x"06537573",
  4392 => x"278d3888",
  4393 => x"15085574",
  4394 => x"782e0981",
  4395 => x"06ea388c",
  4396 => x"150882c8",
  4397 => x"9c0b8405",
  4398 => x"08718c1a",
  4399 => x"0c76881a",
  4400 => x"0c788813",
  4401 => x"0c788c18",
  4402 => x"0c5d5879",
  4403 => x"53807a24",
  4404 => x"83e63872",
  4405 => x"822c8171",
  4406 => x"2b5c537a",
  4407 => x"7c268198",
  4408 => x"387b7b06",
  4409 => x"537282f1",
  4410 => x"3879fc06",
  4411 => x"84055a7a",
  4412 => x"10707d06",
  4413 => x"545b7282",
  4414 => x"e038841a",
  4415 => x"5af13988",
  4416 => x"178c1108",
  4417 => x"58587678",
  4418 => x"2e098106",
  4419 => x"fcc23882",
  4420 => x"1a5afdec",
  4421 => x"39781779",
  4422 => x"81078419",
  4423 => x"0c7082c8",
  4424 => x"b00c7082",
  4425 => x"c8ac0c82",
  4426 => x"c8a40b8c",
  4427 => x"120c8c11",
  4428 => x"0888120c",
  4429 => x"74810784",
  4430 => x"120c7411",
  4431 => x"75710c51",
  4432 => x"537d518b",
  4433 => x"a83f8817",
  4434 => x"54fcac39",
  4435 => x"82c89c0b",
  4436 => x"8405087a",
  4437 => x"545c7980",
  4438 => x"25fef838",
  4439 => x"82da397a",
  4440 => x"097c0670",
  4441 => x"82c89c0b",
  4442 => x"84050c5c",
  4443 => x"7a105b7a",
  4444 => x"7c268538",
  4445 => x"7a85b838",
  4446 => x"82c89c0b",
  4447 => x"88050870",
  4448 => x"841208fc",
  4449 => x"06707c31",
  4450 => x"7c72268f",
  4451 => x"72250757",
  4452 => x"575c5d55",
  4453 => x"72802e80",
  4454 => x"db38797a",
  4455 => x"1682c894",
  4456 => x"081b9011",
  4457 => x"5a55575b",
  4458 => x"82c89008",
  4459 => x"ff2e8838",
  4460 => x"a08f13e0",
  4461 => x"80065776",
  4462 => x"527d51aa",
  4463 => x"f73f8008",
  4464 => x"548008ff",
  4465 => x"2e903880",
  4466 => x"08762782",
  4467 => x"99387482",
  4468 => x"c89c2e82",
  4469 => x"913882c8",
  4470 => x"9c0b8805",
  4471 => x"08558415",
  4472 => x"08fc0670",
  4473 => x"7a317a72",
  4474 => x"268f7225",
  4475 => x"07525553",
  4476 => x"7283e638",
  4477 => x"74798107",
  4478 => x"84170c79",
  4479 => x"167082c8",
  4480 => x"9c0b8805",
  4481 => x"0c758107",
  4482 => x"84120c54",
  4483 => x"7e525789",
  4484 => x"dc3f8817",
  4485 => x"54fae039",
  4486 => x"75832a70",
  4487 => x"54548074",
  4488 => x"24819b38",
  4489 => x"72822c81",
  4490 => x"712b82c8",
  4491 => x"a0080770",
  4492 => x"82c89c0b",
  4493 => x"84050c75",
  4494 => x"10101082",
  4495 => x"c89c0588",
  4496 => x"1108585a",
  4497 => x"5d53778c",
  4498 => x"180c7488",
  4499 => x"180c7688",
  4500 => x"190c768c",
  4501 => x"160cfcf3",
  4502 => x"39797a10",
  4503 => x"101082c8",
  4504 => x"9c057057",
  4505 => x"595d8c15",
  4506 => x"08577675",
  4507 => x"2ea33884",
  4508 => x"1708fc06",
  4509 => x"707a3155",
  4510 => x"56738f24",
  4511 => x"83ca3873",
  4512 => x"80258481",
  4513 => x"388c1708",
  4514 => x"5776752e",
  4515 => x"098106df",
  4516 => x"38881581",
  4517 => x"1b708306",
  4518 => x"555b5572",
  4519 => x"c9387c83",
  4520 => x"06537280",
  4521 => x"2efdb838",
  4522 => x"ff1df819",
  4523 => x"595d8818",
  4524 => x"08782eea",
  4525 => x"38fdb539",
  4526 => x"831a53fc",
  4527 => x"96398314",
  4528 => x"70822c81",
  4529 => x"712b82c8",
  4530 => x"a0080770",
  4531 => x"82c89c0b",
  4532 => x"84050c76",
  4533 => x"10101082",
  4534 => x"c89c0588",
  4535 => x"1108595b",
  4536 => x"5e5153fe",
  4537 => x"e13982c7",
  4538 => x"e0081758",
  4539 => x"8008762e",
  4540 => x"818d3882",
  4541 => x"c89008ff",
  4542 => x"2e83ec38",
  4543 => x"73763118",
  4544 => x"82c7e00c",
  4545 => x"73870670",
  4546 => x"57537280",
  4547 => x"2e883888",
  4548 => x"73317015",
  4549 => x"55567614",
  4550 => x"9fff06a0",
  4551 => x"80713117",
  4552 => x"70547f53",
  4553 => x"5753a88c",
  4554 => x"3f800853",
  4555 => x"8008ff2e",
  4556 => x"81a03882",
  4557 => x"c7e00816",
  4558 => x"7082c7e0",
  4559 => x"0c747582",
  4560 => x"c89c0b88",
  4561 => x"050c7476",
  4562 => x"31187081",
  4563 => x"07515556",
  4564 => x"587b82c8",
  4565 => x"9c2e839c",
  4566 => x"38798f26",
  4567 => x"82cb3881",
  4568 => x"0b84150c",
  4569 => x"841508fc",
  4570 => x"06707a31",
  4571 => x"7a72268f",
  4572 => x"72250752",
  4573 => x"55537280",
  4574 => x"2efcf938",
  4575 => x"80db3980",
  4576 => x"089fff06",
  4577 => x"5372feeb",
  4578 => x"387782c7",
  4579 => x"e00c82c8",
  4580 => x"9c0b8805",
  4581 => x"087b1881",
  4582 => x"0784120c",
  4583 => x"5582c88c",
  4584 => x"08782786",
  4585 => x"387782c8",
  4586 => x"8c0c82c8",
  4587 => x"88087827",
  4588 => x"fcac3877",
  4589 => x"82c8880c",
  4590 => x"841508fc",
  4591 => x"06707a31",
  4592 => x"7a72268f",
  4593 => x"72250752",
  4594 => x"55537280",
  4595 => x"2efca538",
  4596 => x"88398074",
  4597 => x"5456fedb",
  4598 => x"397d5186",
  4599 => x"903f800b",
  4600 => x"800c8f3d",
  4601 => x"0d047353",
  4602 => x"807424a9",
  4603 => x"3872822c",
  4604 => x"81712b82",
  4605 => x"c8a00807",
  4606 => x"7082c89c",
  4607 => x"0b84050c",
  4608 => x"5d53778c",
  4609 => x"180c7488",
  4610 => x"180c7688",
  4611 => x"190c768c",
  4612 => x"160cf9b7",
  4613 => x"39831470",
  4614 => x"822c8171",
  4615 => x"2b82c8a0",
  4616 => x"08077082",
  4617 => x"c89c0b84",
  4618 => x"050c5e51",
  4619 => x"53d4397b",
  4620 => x"7b065372",
  4621 => x"fca33884",
  4622 => x"1a7b105c",
  4623 => x"5af139ff",
  4624 => x"1a811151",
  4625 => x"5af7b939",
  4626 => x"78177981",
  4627 => x"0784190c",
  4628 => x"8c180888",
  4629 => x"1908718c",
  4630 => x"120c8812",
  4631 => x"0c597082",
  4632 => x"c8b00c70",
  4633 => x"82c8ac0c",
  4634 => x"82c8a40b",
  4635 => x"8c120c8c",
  4636 => x"11088812",
  4637 => x"0c748107",
  4638 => x"84120c74",
  4639 => x"1175710c",
  4640 => x"5153f9bd",
  4641 => x"39751784",
  4642 => x"11088107",
  4643 => x"84120c53",
  4644 => x"8c170888",
  4645 => x"1808718c",
  4646 => x"120c8812",
  4647 => x"0c587d51",
  4648 => x"84cb3f88",
  4649 => x"1754f5cf",
  4650 => x"39728415",
  4651 => x"0cf41af8",
  4652 => x"0670841e",
  4653 => x"08810607",
  4654 => x"841e0c70",
  4655 => x"1d545b85",
  4656 => x"0b84140c",
  4657 => x"850b8814",
  4658 => x"0c8f7b27",
  4659 => x"fdcf3888",
  4660 => x"1c527d51",
  4661 => x"e59b3f82",
  4662 => x"c89c0b88",
  4663 => x"050882c7",
  4664 => x"e0085955",
  4665 => x"fdb73977",
  4666 => x"82c7e00c",
  4667 => x"7382c890",
  4668 => x"0cfc9139",
  4669 => x"7284150c",
  4670 => x"fda339fa",
  4671 => x"3d0d7a79",
  4672 => x"028805a7",
  4673 => x"05335652",
  4674 => x"53837327",
  4675 => x"8a387083",
  4676 => x"06527180",
  4677 => x"2ea838ff",
  4678 => x"135372ff",
  4679 => x"2e973870",
  4680 => x"33527372",
  4681 => x"2e913881",
  4682 => x"11ff1454",
  4683 => x"5172ff2e",
  4684 => x"098106eb",
  4685 => x"38805170",
  4686 => x"800c883d",
  4687 => x"0d047072",
  4688 => x"57558351",
  4689 => x"75828029",
  4690 => x"14ff1252",
  4691 => x"56708025",
  4692 => x"f3388373",
  4693 => x"27bf3874",
  4694 => x"08763270",
  4695 => x"09f7fbfd",
  4696 => x"ff120670",
  4697 => x"f8848281",
  4698 => x"80065151",
  4699 => x"5170802e",
  4700 => x"99387451",
  4701 => x"80527033",
  4702 => x"5773772e",
  4703 => x"ffb93881",
  4704 => x"11811353",
  4705 => x"51837227",
  4706 => x"ed38fc13",
  4707 => x"84165653",
  4708 => x"728326c3",
  4709 => x"387451fe",
  4710 => x"fe39fa3d",
  4711 => x"0d787a7c",
  4712 => x"72727257",
  4713 => x"57575956",
  4714 => x"56747627",
  4715 => x"b2387615",
  4716 => x"51757127",
  4717 => x"aa387077",
  4718 => x"17ff1454",
  4719 => x"555371ff",
  4720 => x"2e9638ff",
  4721 => x"14ff1454",
  4722 => x"54723374",
  4723 => x"34ff1252",
  4724 => x"71ff2e09",
  4725 => x"8106ec38",
  4726 => x"75800c88",
  4727 => x"3d0d0476",
  4728 => x"8f269738",
  4729 => x"ff125271",
  4730 => x"ff2eed38",
  4731 => x"72708105",
  4732 => x"54337470",
  4733 => x"81055634",
  4734 => x"eb397476",
  4735 => x"07830651",
  4736 => x"70e23875",
  4737 => x"75545172",
  4738 => x"70840554",
  4739 => x"08717084",
  4740 => x"05530c72",
  4741 => x"70840554",
  4742 => x"08717084",
  4743 => x"05530c72",
  4744 => x"70840554",
  4745 => x"08717084",
  4746 => x"05530c72",
  4747 => x"70840554",
  4748 => x"08717084",
  4749 => x"05530cf0",
  4750 => x"1252718f",
  4751 => x"26c93883",
  4752 => x"72279538",
  4753 => x"72708405",
  4754 => x"54087170",
  4755 => x"8405530c",
  4756 => x"fc125271",
  4757 => x"8326ed38",
  4758 => x"7054ff88",
  4759 => x"39fc3d0d",
  4760 => x"76797102",
  4761 => x"8c059f05",
  4762 => x"33575553",
  4763 => x"55837227",
  4764 => x"8a387483",
  4765 => x"06517080",
  4766 => x"2ea238ff",
  4767 => x"125271ff",
  4768 => x"2e933873",
  4769 => x"73708105",
  4770 => x"5534ff12",
  4771 => x"5271ff2e",
  4772 => x"098106ef",
  4773 => x"3874800c",
  4774 => x"863d0d04",
  4775 => x"7474882b",
  4776 => x"75077071",
  4777 => x"902b0751",
  4778 => x"54518f72",
  4779 => x"27a53872",
  4780 => x"71708405",
  4781 => x"530c7271",
  4782 => x"70840553",
  4783 => x"0c727170",
  4784 => x"8405530c",
  4785 => x"72717084",
  4786 => x"05530cf0",
  4787 => x"1252718f",
  4788 => x"26dd3883",
  4789 => x"72279038",
  4790 => x"72717084",
  4791 => x"05530cfc",
  4792 => x"12527183",
  4793 => x"26f23870",
  4794 => x"53ff9039",
  4795 => x"0404f93d",
  4796 => x"0d797b80",
  4797 => x"cc120856",
  4798 => x"58567380",
  4799 => x"2ea53876",
  4800 => x"10101470",
  4801 => x"08555573",
  4802 => x"802eb538",
  4803 => x"7308750c",
  4804 => x"800b9015",
  4805 => x"0c800b8c",
  4806 => x"150c7355",
  4807 => x"74800c89",
  4808 => x"3d0d0490",
  4809 => x"53845275",
  4810 => x"51a5f63f",
  4811 => x"800880cc",
  4812 => x"170c8008",
  4813 => x"55800880",
  4814 => x"2ee23880",
  4815 => x"0854c039",
  4816 => x"81772b70",
  4817 => x"10109405",
  4818 => x"54588152",
  4819 => x"7551a5d1",
  4820 => x"3f800880",
  4821 => x"08565480",
  4822 => x"08802ec0",
  4823 => x"38768008",
  4824 => x"84050c77",
  4825 => x"80088805",
  4826 => x"0c800b90",
  4827 => x"150c800b",
  4828 => x"8c150c73",
  4829 => x"55ffa539",
  4830 => x"ff3d0d74",
  4831 => x"5271802e",
  4832 => x"95387384",
  4833 => x"13081010",
  4834 => x"80cc1208",
  4835 => x"05700874",
  4836 => x"0c73710c",
  4837 => x"5151833d",
  4838 => x"0d04f53d",
  4839 => x"0d7d7f61",
  4840 => x"63901308",
  4841 => x"94145b5d",
  4842 => x"5b5c5c5c",
  4843 => x"80578216",
  4844 => x"227a7129",
  4845 => x"1977227c",
  4846 => x"71297290",
  4847 => x"2a057090",
  4848 => x"2a7383ff",
  4849 => x"ff067284",
  4850 => x"80802905",
  4851 => x"7b708405",
  4852 => x"5d0c811c",
  4853 => x"5c52535a",
  4854 => x"55557877",
  4855 => x"24d03877",
  4856 => x"802e9638",
  4857 => x"78881c08",
  4858 => x"25963878",
  4859 => x"10101b78",
  4860 => x"94120c54",
  4861 => x"8119901c",
  4862 => x"0c7a800c",
  4863 => x"8d3d0d04",
  4864 => x"841b0881",
  4865 => x"05527b51",
  4866 => x"fde43f80",
  4867 => x"08901c08",
  4868 => x"10108805",
  4869 => x"548c1c53",
  4870 => x"80088c05",
  4871 => x"5254fef9",
  4872 => x"ee3f7a52",
  4873 => x"7b51fed0",
  4874 => x"3f737910",
  4875 => x"10117994",
  4876 => x"120c5581",
  4877 => x"1a90120c",
  4878 => x"5bffbe39",
  4879 => x"f63d0d7c",
  4880 => x"7e60625e",
  4881 => x"5c595989",
  4882 => x"52881b51",
  4883 => x"fef5903f",
  4884 => x"80085780",
  4885 => x"56815574",
  4886 => x"77258c38",
  4887 => x"74108117",
  4888 => x"57557675",
  4889 => x"24f63875",
  4890 => x"527851fd",
  4891 => x"813f8008",
  4892 => x"61800894",
  4893 => x"050c5681",
  4894 => x"0b800890",
  4895 => x"050c8957",
  4896 => x"767a2580",
  4897 => x"cf387618",
  4898 => x"58777081",
  4899 => x"055933d0",
  4900 => x"05548a53",
  4901 => x"75527851",
  4902 => x"fe803f80",
  4903 => x"08811858",
  4904 => x"56797724",
  4905 => x"e4388118",
  4906 => x"58767b25",
  4907 => x"a0387a77",
  4908 => x"31577770",
  4909 => x"81055933",
  4910 => x"d005548a",
  4911 => x"53755278",
  4912 => x"51fdd73f",
  4913 => x"8008ff18",
  4914 => x"585676e6",
  4915 => x"3875800c",
  4916 => x"8c3d0d04",
  4917 => x"8a1858d1",
  4918 => x"39fe3d0d",
  4919 => x"74528072",
  4920 => x"fc808006",
  4921 => x"52537073",
  4922 => x"2e098106",
  4923 => x"87389072",
  4924 => x"712b5353",
  4925 => x"7181ff0a",
  4926 => x"06517088",
  4927 => x"38881372",
  4928 => x"882b5353",
  4929 => x"718f0a06",
  4930 => x"51708838",
  4931 => x"84137284",
  4932 => x"2b535371",
  4933 => x"830a0651",
  4934 => x"70883882",
  4935 => x"1372822b",
  4936 => x"53538072",
  4937 => x"24933881",
  4938 => x"13729e2a",
  4939 => x"70810651",
  4940 => x"5253a052",
  4941 => x"70802e83",
  4942 => x"38725271",
  4943 => x"800c843d",
  4944 => x"0d04fc3d",
  4945 => x"0d767008",
  4946 => x"70870653",
  4947 => x"53557080",
  4948 => x"2eaa3871",
  4949 => x"81065180",
  4950 => x"5370732e",
  4951 => x"09810695",
  4952 => x"38710a10",
  4953 => x"0a708106",
  4954 => x"52537080",
  4955 => x"2e80f038",
  4956 => x"72750c81",
  4957 => x"5372800c",
  4958 => x"863d0d04",
  4959 => x"707283ff",
  4960 => x"ff065254",
  4961 => x"70802e80",
  4962 => x"cd387181",
  4963 => x"ff065170",
  4964 => x"88388814",
  4965 => x"72882a53",
  4966 => x"54718f06",
  4967 => x"51708838",
  4968 => x"84147284",
  4969 => x"2a535471",
  4970 => x"83065170",
  4971 => x"88388214",
  4972 => x"72822a53",
  4973 => x"54718106",
  4974 => x"51709138",
  4975 => x"8114720a",
  4976 => x"100a5354",
  4977 => x"a0537180",
  4978 => x"2effaa38",
  4979 => x"71750c73",
  4980 => x"800c863d",
  4981 => x"0d049072",
  4982 => x"712a5354",
  4983 => x"ffac3971",
  4984 => x"822a750c",
  4985 => x"820b800c",
  4986 => x"863d0d04",
  4987 => x"ff3d0d81",
  4988 => x"527351f9",
  4989 => x"f93f7480",
  4990 => x"0894050c",
  4991 => x"810b8008",
  4992 => x"90050c83",
  4993 => x"3d0d04ee",
  4994 => x"3d0d6567",
  4995 => x"90120890",
  4996 => x"12085856",
  4997 => x"57537375",
  4998 => x"258d3872",
  4999 => x"76717790",
  5000 => x"14085957",
  5001 => x"58544274",
  5002 => x"14708815",
  5003 => x"08248415",
  5004 => x"08055365",
  5005 => x"525ef9b6",
  5006 => x"3f800880",
  5007 => x"08940570",
  5008 => x"60822b72",
  5009 => x"11434659",
  5010 => x"41427f7f",
  5011 => x"278d3880",
  5012 => x"77708405",
  5013 => x"590c7e77",
  5014 => x"26f53894",
  5015 => x"13741010",
  5016 => x"11941877",
  5017 => x"10101163",
  5018 => x"41445d5d",
  5019 => x"5f7a6127",
  5020 => x"81b8387a",
  5021 => x"087083ff",
  5022 => x"ff065953",
  5023 => x"77802e80",
  5024 => x"c7387e7d",
  5025 => x"5757805a",
  5026 => x"76708405",
  5027 => x"58087083",
  5028 => x"ffff0682",
  5029 => x"1822717b",
  5030 => x"29057c11",
  5031 => x"73902a7c",
  5032 => x"297a225e",
  5033 => x"7d057190",
  5034 => x"2a057090",
  5035 => x"2a5f5951",
  5036 => x"51545474",
  5037 => x"76237282",
  5038 => x"17238416",
  5039 => x"567b7726",
  5040 => x"c7387976",
  5041 => x"0c7a0853",
  5042 => x"72902a58",
  5043 => x"77802e80",
  5044 => x"cd387e7d",
  5045 => x"5757807d",
  5046 => x"08705b56",
  5047 => x"5a767084",
  5048 => x"05580870",
  5049 => x"83ffff06",
  5050 => x"707a297b",
  5051 => x"902a057c",
  5052 => x"11515154",
  5053 => x"54727623",
  5054 => x"74821723",
  5055 => x"84167490",
  5056 => x"2a792971",
  5057 => x"08821322",
  5058 => x"5d5b7b05",
  5059 => x"74902a05",
  5060 => x"70902a5c",
  5061 => x"56567b77",
  5062 => x"26c33874",
  5063 => x"760c841b",
  5064 => x"841e5e5b",
  5065 => x"607b26fe",
  5066 => x"ca386260",
  5067 => x"0556807e",
  5068 => x"259038fc",
  5069 => x"16567508",
  5070 => x"8938ff1e",
  5071 => x"5e7d8024",
  5072 => x"f2387d62",
  5073 => x"90050c61",
  5074 => x"800c943d",
  5075 => x"0d04f73d",
  5076 => x"0d7b7d7f",
  5077 => x"70830658",
  5078 => x"585a5a74",
  5079 => x"80dd3875",
  5080 => x"822c5675",
  5081 => x"802eb638",
  5082 => x"80c81a08",
  5083 => x"70565776",
  5084 => x"802e80f8",
  5085 => x"38758106",
  5086 => x"5574a938",
  5087 => x"75812c56",
  5088 => x"75802e99",
  5089 => x"38760870",
  5090 => x"59557480",
  5091 => x"2e80c638",
  5092 => x"74577581",
  5093 => x"06557480",
  5094 => x"2ee23888",
  5095 => x"3978800c",
  5096 => x"8b3d0d04",
  5097 => x"76537852",
  5098 => x"7951fcdb",
  5099 => x"3f800879",
  5100 => x"537a5255",
  5101 => x"f7c23f74",
  5102 => x"59c23980",
  5103 => x"54741010",
  5104 => x"82bff005",
  5105 => x"70085455",
  5106 => x"78527951",
  5107 => x"f7cc3f80",
  5108 => x"0859ff8b",
  5109 => x"39765376",
  5110 => x"527951fc",
  5111 => x"aa3f8008",
  5112 => x"770c8008",
  5113 => x"7880080c",
  5114 => x"57ffa739",
  5115 => x"84f15279",
  5116 => x"51fbf93f",
  5117 => x"800880c8",
  5118 => x"1b0c8008",
  5119 => x"7580080c",
  5120 => x"76810656",
  5121 => x"5774802e",
  5122 => x"fef238ff",
  5123 => x"9739f53d",
  5124 => x"0d7d7f61",
  5125 => x"70852c84",
  5126 => x"13089014",
  5127 => x"08128105",
  5128 => x"88150859",
  5129 => x"5e59595a",
  5130 => x"5c5c7279",
  5131 => x"258c3881",
  5132 => x"15731054",
  5133 => x"55787324",
  5134 => x"f6387452",
  5135 => x"7b51f5ae",
  5136 => x"3f800880",
  5137 => x"08940555",
  5138 => x"5a807625",
  5139 => x"90387553",
  5140 => x"80747084",
  5141 => x"05560cff",
  5142 => x"135372f4",
  5143 => x"38941b90",
  5144 => x"1c081010",
  5145 => x"11799f06",
  5146 => x"5a585377",
  5147 => x"802ebf38",
  5148 => x"a0783155",
  5149 => x"80567208",
  5150 => x"782b7607",
  5151 => x"74708405",
  5152 => x"560c7270",
  5153 => x"84055408",
  5154 => x"752a5676",
  5155 => x"7326e738",
  5156 => x"75740c75",
  5157 => x"802e8438",
  5158 => x"811959ff",
  5159 => x"19901b0c",
  5160 => x"7a527b51",
  5161 => x"f5d23f79",
  5162 => x"800c8d3d",
  5163 => x"0d047270",
  5164 => x"84055408",
  5165 => x"74708405",
  5166 => x"560c7277",
  5167 => x"27dd3872",
  5168 => x"70840554",
  5169 => x"08747084",
  5170 => x"05560c76",
  5171 => x"7326df38",
  5172 => x"ca39fb3d",
  5173 => x"0d777990",
  5174 => x"11089013",
  5175 => x"08713170",
  5176 => x"56545557",
  5177 => x"5470ab38",
  5178 => x"94147382",
  5179 => x"2b711171",
  5180 => x"19940552",
  5181 => x"545255fc",
  5182 => x"12fc1271",
  5183 => x"08710856",
  5184 => x"56525273",
  5185 => x"732e0981",
  5186 => x"068f3871",
  5187 => x"7526e838",
  5188 => x"80527180",
  5189 => x"0c873d0d",
  5190 => x"04ff5172",
  5191 => x"74268338",
  5192 => x"81517080",
  5193 => x"0c873d0d",
  5194 => x"04f33d0d",
  5195 => x"7f616370",
  5196 => x"55715457",
  5197 => x"5456ff9a",
  5198 => x"3f800854",
  5199 => x"8008802e",
  5200 => x"81c63880",
  5201 => x"54738008",
  5202 => x"2481dc38",
  5203 => x"84130852",
  5204 => x"7551f39a",
  5205 => x"3f800874",
  5206 => x"80088c05",
  5207 => x"0c901408",
  5208 => x"94157110",
  5209 => x"10119419",
  5210 => x"901a0810",
  5211 => x"10118008",
  5212 => x"94055d41",
  5213 => x"5d415a5c",
  5214 => x"5d805a77",
  5215 => x"70840559",
  5216 => x"087083ff",
  5217 => x"ff067a70",
  5218 => x"84055c08",
  5219 => x"7083ffff",
  5220 => x"06727131",
  5221 => x"1e74902a",
  5222 => x"73902a31",
  5223 => x"71902c11",
  5224 => x"70902c41",
  5225 => x"51555156",
  5226 => x"57575473",
  5227 => x"77237282",
  5228 => x"18238417",
  5229 => x"577b7926",
  5230 => x"c238777e",
  5231 => x"27ac3877",
  5232 => x"70840559",
  5233 => x"087083ff",
  5234 => x"ff067b11",
  5235 => x"70902c73",
  5236 => x"902a0570",
  5237 => x"902c5e53",
  5238 => x"51545473",
  5239 => x"77237282",
  5240 => x"18238417",
  5241 => x"577d7826",
  5242 => x"d638fc17",
  5243 => x"5776088d",
  5244 => x"38ff1bfc",
  5245 => x"18585b76",
  5246 => x"08802ef5",
  5247 => x"387a901e",
  5248 => x"0c7c800c",
  5249 => x"8f3d0d04",
  5250 => x"80085275",
  5251 => x"51f1df3f",
  5252 => x"80085d81",
  5253 => x"0b800890",
  5254 => x"050c7380",
  5255 => x"0894050c",
  5256 => x"7c800c8f",
  5257 => x"3d0d0472",
  5258 => x"75545581",
  5259 => x"0b841408",
  5260 => x"53765254",
  5261 => x"f1b83f80",
  5262 => x"08748008",
  5263 => x"8c050c90",
  5264 => x"14089415",
  5265 => x"71101011",
  5266 => x"9419901a",
  5267 => x"08101011",
  5268 => x"80089405",
  5269 => x"5d415d41",
  5270 => x"5a5c5d80",
  5271 => x"5afe9c39",
  5272 => x"fa3d0d78",
  5273 => x"7a7c5457",
  5274 => x"7258769f",
  5275 => x"fe0a0686",
  5276 => x"bf0a0553",
  5277 => x"53807225",
  5278 => x"95387154",
  5279 => x"80557375",
  5280 => x"53730c71",
  5281 => x"84140c72",
  5282 => x"800c883d",
  5283 => x"0d047130",
  5284 => x"70942c53",
  5285 => x"51937225",
  5286 => x"a7388054",
  5287 => x"ec129f71",
  5288 => x"3181712b",
  5289 => x"5152529e",
  5290 => x"72258338",
  5291 => x"81517055",
  5292 => x"73755373",
  5293 => x"0c718414",
  5294 => x"0c72800c",
  5295 => x"883d0d04",
  5296 => x"a0808072",
  5297 => x"2c548055",
  5298 => x"ffb439f6",
  5299 => x"3d0d7c7e",
  5300 => x"94119012",
  5301 => x"08101011",
  5302 => x"fc117008",
  5303 => x"70575a51",
  5304 => x"57585359",
  5305 => x"f3f33f80",
  5306 => x"087fa00b",
  5307 => x"80083171",
  5308 => x"0c53538a",
  5309 => x"0b800825",
  5310 => x"80e83880",
  5311 => x"57737626",
  5312 => x"bd38f513",
  5313 => x"5372802e",
  5314 => x"80c038a0",
  5315 => x"73317574",
  5316 => x"2b78722a",
  5317 => x"079ffc0a",
  5318 => x"075b5880",
  5319 => x"55757427",
  5320 => x"8538fc14",
  5321 => x"08557673",
  5322 => x"2b75792a",
  5323 => x"075b797b",
  5324 => x"54790c72",
  5325 => x"841a0c78",
  5326 => x"800c8c3d",
  5327 => x"0d04fc14",
  5328 => x"7008f515",
  5329 => x"55585472",
  5330 => x"c238749f",
  5331 => x"fc0a075a",
  5332 => x"765b797b",
  5333 => x"54790c72",
  5334 => x"841a0c78",
  5335 => x"800c8c3d",
  5336 => x"0d048b0b",
  5337 => x"80083175",
  5338 => x"712a9ffc",
  5339 => x"0a075b57",
  5340 => x"80587574",
  5341 => x"278538fc",
  5342 => x"14085895",
  5343 => x"1375712b",
  5344 => x"79792a07",
  5345 => x"5c52797b",
  5346 => x"54790c72",
  5347 => x"841a0c78",
  5348 => x"800c8c3d",
  5349 => x"0d04f33d",
  5350 => x"0d626462",
  5351 => x"64575f75",
  5352 => x"405b5981",
  5353 => x"527f51ee",
  5354 => x"c53f8008",
  5355 => x"80089405",
  5356 => x"7e70bfff",
  5357 => x"ff06705f",
  5358 => x"71fe0a06",
  5359 => x"70427094",
  5360 => x"2a5b5257",
  5361 => x"55595775",
  5362 => x"802e8738",
  5363 => x"7390800a",
  5364 => x"075b7d53",
  5365 => x"72802e80",
  5366 => x"d638725c",
  5367 => x"8f3df405",
  5368 => x"51f2df3f",
  5369 => x"80085580",
  5370 => x"08802e80",
  5371 => x"ff38a00b",
  5372 => x"8008317b",
  5373 => x"712b7d07",
  5374 => x"790c537a",
  5375 => x"80082a5b",
  5376 => x"7a70841a",
  5377 => x"0c703070",
  5378 => x"72078025",
  5379 => x"82713170",
  5380 => x"901c0c51",
  5381 => x"51545475",
  5382 => x"802eaf38",
  5383 => x"7416f7cd",
  5384 => x"05790cb5",
  5385 => x"75317a0c",
  5386 => x"76800c8f",
  5387 => x"3d0d048f",
  5388 => x"3df00551",
  5389 => x"f28c3f7a",
  5390 => x"780c810b",
  5391 => x"90180c81",
  5392 => x"0b8008a0",
  5393 => x"05565375",
  5394 => x"d338f7ce",
  5395 => x"15790c72",
  5396 => x"852b7310",
  5397 => x"1019fc11",
  5398 => x"08535454",
  5399 => x"f0fb3f73",
  5400 => x"8008317a",
  5401 => x"0c76800c",
  5402 => x"8f3d0d04",
  5403 => x"7b780c7a",
  5404 => x"70841a0c",
  5405 => x"70307072",
  5406 => x"07802582",
  5407 => x"71317090",
  5408 => x"1c0c5151",
  5409 => x"5454ff8f",
  5410 => x"39f03d0d",
  5411 => x"62646695",
  5412 => x"3de41157",
  5413 => x"7256f805",
  5414 => x"54585858",
  5415 => x"fcad3f92",
  5416 => x"3de01154",
  5417 => x"7653f005",
  5418 => x"51fca03f",
  5419 => x"90170890",
  5420 => x"17083185",
  5421 => x"2b7b7b31",
  5422 => x"11515680",
  5423 => x"7625ae38",
  5424 => x"7590800a",
  5425 => x"29600540",
  5426 => x"7d7f5854",
  5427 => x"76557f61",
  5428 => x"58527653",
  5429 => x"923de805",
  5430 => x"5180cbb7",
  5431 => x"3f7b7d58",
  5432 => x"780c7684",
  5433 => x"190c7780",
  5434 => x"0c923d0d",
  5435 => x"04753070",
  5436 => x"90800a29",
  5437 => x"1f5f567d",
  5438 => x"7f585476",
  5439 => x"557f6158",
  5440 => x"52765392",
  5441 => x"3de80551",
  5442 => x"80cb883f",
  5443 => x"7b7d5878",
  5444 => x"0c768419",
  5445 => x"0c77800c",
  5446 => x"923d0d04",
  5447 => x"f33d0d7f",
  5448 => x"61575c9f",
  5449 => x"fc0a5780",
  5450 => x"58759724",
  5451 => x"9b387510",
  5452 => x"101082be",
  5453 => x"ac058411",
  5454 => x"0871087e",
  5455 => x"0c841e0c",
  5456 => x"7c800c56",
  5457 => x"8f3d0d04",
  5458 => x"807625a4",
  5459 => x"388d3d5b",
  5460 => x"80c8820a",
  5461 => x"59805a78",
  5462 => x"54795576",
  5463 => x"5277537a",
  5464 => x"51ada13f",
  5465 => x"7c7eff18",
  5466 => x"58595775",
  5467 => x"8024e838",
  5468 => x"767c0c77",
  5469 => x"841d0c7b",
  5470 => x"800c8f3d",
  5471 => x"0d04ef3d",
  5472 => x"0d636567",
  5473 => x"405d427b",
  5474 => x"802e84fa",
  5475 => x"386151ea",
  5476 => x"db3ff81c",
  5477 => x"70841208",
  5478 => x"70fc0670",
  5479 => x"628b0570",
  5480 => x"f8064159",
  5481 => x"455b5c41",
  5482 => x"57967427",
  5483 => x"82c33880",
  5484 => x"7b247e7c",
  5485 => x"26075980",
  5486 => x"5478742e",
  5487 => x"09810682",
  5488 => x"a938777b",
  5489 => x"2581fc38",
  5490 => x"771782c8",
  5491 => x"9c0b8805",
  5492 => x"085e567c",
  5493 => x"762e84bd",
  5494 => x"38841608",
  5495 => x"70fe0617",
  5496 => x"84110881",
  5497 => x"06515555",
  5498 => x"73828b38",
  5499 => x"74fc0659",
  5500 => x"7c762e84",
  5501 => x"de387719",
  5502 => x"5f7e7b25",
  5503 => x"81fd3879",
  5504 => x"81065473",
  5505 => x"82bf3876",
  5506 => x"77083184",
  5507 => x"1108fc06",
  5508 => x"565a7580",
  5509 => x"2e91387c",
  5510 => x"762e84eb",
  5511 => x"38741918",
  5512 => x"59787b25",
  5513 => x"848a3879",
  5514 => x"802e8299",
  5515 => x"38771556",
  5516 => x"7a762482",
  5517 => x"90388c1a",
  5518 => x"08881b08",
  5519 => x"718c120c",
  5520 => x"88120c55",
  5521 => x"79765957",
  5522 => x"881761fc",
  5523 => x"05575975",
  5524 => x"a42685f0",
  5525 => x"387b7955",
  5526 => x"55937627",
  5527 => x"80c9387b",
  5528 => x"7084055d",
  5529 => x"087c5679",
  5530 => x"0c747084",
  5531 => x"0556088c",
  5532 => x"180c9017",
  5533 => x"549b7627",
  5534 => x"ae387470",
  5535 => x"84055608",
  5536 => x"740c7470",
  5537 => x"84055608",
  5538 => x"94180c98",
  5539 => x"1754a376",
  5540 => x"27953874",
  5541 => x"70840556",
  5542 => x"08740c74",
  5543 => x"70840556",
  5544 => x"089c180c",
  5545 => x"a0175474",
  5546 => x"70840556",
  5547 => x"08747084",
  5548 => x"05560c74",
  5549 => x"70840556",
  5550 => x"08747084",
  5551 => x"05560c74",
  5552 => x"08740c77",
  5553 => x"7b315675",
  5554 => x"8f2680c9",
  5555 => x"38841708",
  5556 => x"81067807",
  5557 => x"84180c77",
  5558 => x"17841108",
  5559 => x"81078412",
  5560 => x"0c546151",
  5561 => x"e8873f88",
  5562 => x"17547380",
  5563 => x"0c933d0d",
  5564 => x"04905bfd",
  5565 => x"ba397856",
  5566 => x"fe85398c",
  5567 => x"16088817",
  5568 => x"08718c12",
  5569 => x"0c88120c",
  5570 => x"557e707c",
  5571 => x"3157588f",
  5572 => x"7627ffb9",
  5573 => x"387a1784",
  5574 => x"18088106",
  5575 => x"7c078419",
  5576 => x"0c768107",
  5577 => x"84120c76",
  5578 => x"11841108",
  5579 => x"81078412",
  5580 => x"0c558805",
  5581 => x"526151c8",
  5582 => x"b83f6151",
  5583 => x"e7af3f88",
  5584 => x"1754ffa6",
  5585 => x"397d5261",
  5586 => x"51d7ba3f",
  5587 => x"80085980",
  5588 => x"08802e81",
  5589 => x"a3388008",
  5590 => x"f8056084",
  5591 => x"0508fe06",
  5592 => x"61055557",
  5593 => x"76742e83",
  5594 => x"e838fc18",
  5595 => x"5675a426",
  5596 => x"81aa387b",
  5597 => x"80085555",
  5598 => x"93762780",
  5599 => x"d8387470",
  5600 => x"84055608",
  5601 => x"80087084",
  5602 => x"05800c0c",
  5603 => x"80087570",
  5604 => x"84055708",
  5605 => x"71708405",
  5606 => x"530c549b",
  5607 => x"7627b638",
  5608 => x"74708405",
  5609 => x"56087470",
  5610 => x"8405560c",
  5611 => x"74708405",
  5612 => x"56087470",
  5613 => x"8405560c",
  5614 => x"a3762799",
  5615 => x"38747084",
  5616 => x"05560874",
  5617 => x"70840556",
  5618 => x"0c747084",
  5619 => x"05560874",
  5620 => x"70840556",
  5621 => x"0c747084",
  5622 => x"05560874",
  5623 => x"70840556",
  5624 => x"0c747084",
  5625 => x"05560874",
  5626 => x"70840556",
  5627 => x"0c740874",
  5628 => x"0c7b5261",
  5629 => x"51c6fa3f",
  5630 => x"6151e5f1",
  5631 => x"3f785473",
  5632 => x"800c933d",
  5633 => x"0d047d52",
  5634 => x"6151d5f9",
  5635 => x"3f800880",
  5636 => x"0c933d0d",
  5637 => x"04841608",
  5638 => x"55fbd139",
  5639 => x"75537b52",
  5640 => x"800851fe",
  5641 => x"e1e93f7b",
  5642 => x"526151c6",
  5643 => x"c43fc939",
  5644 => x"8c160888",
  5645 => x"1708718c",
  5646 => x"120c8812",
  5647 => x"0c558c1a",
  5648 => x"08881b08",
  5649 => x"718c120c",
  5650 => x"88120c55",
  5651 => x"79795957",
  5652 => x"fbf63977",
  5653 => x"19901c55",
  5654 => x"55737524",
  5655 => x"fba1387a",
  5656 => x"177082c8",
  5657 => x"9c0b8805",
  5658 => x"0c757c31",
  5659 => x"81078412",
  5660 => x"0c5d8417",
  5661 => x"0881067b",
  5662 => x"0784180c",
  5663 => x"6151e4ed",
  5664 => x"3f881754",
  5665 => x"fce43974",
  5666 => x"1918901c",
  5667 => x"555d737d",
  5668 => x"24fb9438",
  5669 => x"8c1a0888",
  5670 => x"1b08718c",
  5671 => x"120c8812",
  5672 => x"0c55881a",
  5673 => x"61fc0557",
  5674 => x"5975a426",
  5675 => x"81af387b",
  5676 => x"79555593",
  5677 => x"762780c9",
  5678 => x"387b7084",
  5679 => x"055d087c",
  5680 => x"56790c74",
  5681 => x"70840556",
  5682 => x"088c1b0c",
  5683 => x"901a549b",
  5684 => x"7627ae38",
  5685 => x"74708405",
  5686 => x"5608740c",
  5687 => x"74708405",
  5688 => x"5608941b",
  5689 => x"0c981a54",
  5690 => x"a3762795",
  5691 => x"38747084",
  5692 => x"05560874",
  5693 => x"0c747084",
  5694 => x"0556089c",
  5695 => x"1b0ca01a",
  5696 => x"54747084",
  5697 => x"05560874",
  5698 => x"70840556",
  5699 => x"0c747084",
  5700 => x"05560874",
  5701 => x"70840556",
  5702 => x"0c740874",
  5703 => x"0c7a1a70",
  5704 => x"82c89c0b",
  5705 => x"88050c7d",
  5706 => x"7c318107",
  5707 => x"84120c54",
  5708 => x"841a0881",
  5709 => x"067b0784",
  5710 => x"1b0c6151",
  5711 => x"e3af3f78",
  5712 => x"54fdbc39",
  5713 => x"75537b52",
  5714 => x"7851fedf",
  5715 => x"c23ffaf3",
  5716 => x"39841708",
  5717 => x"fc061860",
  5718 => x"5858fae7",
  5719 => x"3975537b",
  5720 => x"527851fe",
  5721 => x"dfa93f7a",
  5722 => x"1a7082c8",
  5723 => x"9c0b8805",
  5724 => x"0c7d7c31",
  5725 => x"81078412",
  5726 => x"0c54841a",
  5727 => x"0881067b",
  5728 => x"07841b0c",
  5729 => x"ffb439fd",
  5730 => x"3d0d758c",
  5731 => x"11228906",
  5732 => x"53548053",
  5733 => x"71892e88",
  5734 => x"3872800c",
  5735 => x"853d0d04",
  5736 => x"7351ffbc",
  5737 => x"ff3f8008",
  5738 => x"800c853d",
  5739 => x"0d04f93d",
  5740 => x"0d7982c0",
  5741 => x"c0085556",
  5742 => x"b8140880",
  5743 => x"2e81e038",
  5744 => x"800b8c17",
  5745 => x"227083ff",
  5746 => x"ff067085",
  5747 => x"2a708106",
  5748 => x"51575758",
  5749 => x"5873782e",
  5750 => x"09810682",
  5751 => x"a5387482",
  5752 => x"2a813270",
  5753 => x"81065154",
  5754 => x"73802e80",
  5755 => x"f3387784",
  5756 => x"170c7484",
  5757 => x"2a813270",
  5758 => x"81065154",
  5759 => x"ff587380",
  5760 => x"d8387483",
  5761 => x"2a708106",
  5762 => x"51547381",
  5763 => x"c9387684",
  5764 => x"0754738c",
  5765 => x"17239016",
  5766 => x"08802e81",
  5767 => x"9a388c16",
  5768 => x"22830654",
  5769 => x"73818138",
  5770 => x"90160876",
  5771 => x"0c941608",
  5772 => x"53750852",
  5773 => x"9c160851",
  5774 => x"a0160854",
  5775 => x"732d8c16",
  5776 => x"2283bfff",
  5777 => x"0654800b",
  5778 => x"80082581",
  5779 => x"c2388008",
  5780 => x"84170c73",
  5781 => x"8c172380",
  5782 => x"5877800c",
  5783 => x"893d0d04",
  5784 => x"b0160855",
  5785 => x"74802e80",
  5786 => x"e13880c0",
  5787 => x"16547474",
  5788 => x"2e8f3877",
  5789 => x"84170c74",
  5790 => x"5282c0c0",
  5791 => x"0851c1f1",
  5792 => x"3f77b017",
  5793 => x"0cbc1608",
  5794 => x"7084180c",
  5795 => x"5473802e",
  5796 => x"ff8438b8",
  5797 => x"1608760c",
  5798 => x"77800c89",
  5799 => x"3d0d0473",
  5800 => x"51ffbde3",
  5801 => x"3ffe9939",
  5802 => x"81b38752",
  5803 => x"82c0c008",
  5804 => x"51cbfb3f",
  5805 => x"fef23975",
  5806 => x"51cea53f",
  5807 => x"8c162283",
  5808 => x"06547380",
  5809 => x"2efee138",
  5810 => x"df397784",
  5811 => x"170c9016",
  5812 => x"08fecb38",
  5813 => x"e2397551",
  5814 => x"ffbac93f",
  5815 => x"8008fef9",
  5816 => x"388c1622",
  5817 => x"83fff706",
  5818 => x"54738c17",
  5819 => x"23800888",
  5820 => x"170c8008",
  5821 => x"98170c73",
  5822 => x"84075473",
  5823 => x"8c1723fe",
  5824 => x"95397784",
  5825 => x"170cff58",
  5826 => x"77800c89",
  5827 => x"3d0d0480",
  5828 => x"08923880",
  5829 => x"0884170c",
  5830 => x"73a00754",
  5831 => x"738c1723",
  5832 => x"ff58e539",
  5833 => x"800b8417",
  5834 => x"0c7380c0",
  5835 => x"0754738c",
  5836 => x"1723ed39",
  5837 => x"fd3d0d80",
  5838 => x"0b82d0d4",
  5839 => x"0c765188",
  5840 => x"ca3f8008",
  5841 => x"538008ff",
  5842 => x"2e883872",
  5843 => x"800c853d",
  5844 => x"0d0482d0",
  5845 => x"d4085473",
  5846 => x"802ef038",
  5847 => x"7574710c",
  5848 => x"5272800c",
  5849 => x"853d0d04",
  5850 => x"fd3d0d75",
  5851 => x"77535371",
  5852 => x"54733070",
  5853 => x"75079f2a",
  5854 => x"7075fe0a",
  5855 => x"06079081",
  5856 => x"0a119ffe",
  5857 => x"0a723107",
  5858 => x"709f2a81",
  5859 => x"7131800c",
  5860 => x"51515151",
  5861 => x"51853d0d",
  5862 => x"04fd3d0d",
  5863 => x"75775353",
  5864 => x"71547330",
  5865 => x"7075079f",
  5866 => x"2a7075fe",
  5867 => x"0a06079f",
  5868 => x"fe0a7131",
  5869 => x"9f2a800c",
  5870 => x"51515185",
  5871 => x"3d0d04f9",
  5872 => x"3d0d797c",
  5873 => x"557b548e",
  5874 => x"11227090",
  5875 => x"2b70902c",
  5876 => x"555782c0",
  5877 => x"c0085358",
  5878 => x"5686f83f",
  5879 => x"80085780",
  5880 => x"0b800824",
  5881 => x"933880d0",
  5882 => x"16088008",
  5883 => x"0580d017",
  5884 => x"0c76800c",
  5885 => x"893d0d04",
  5886 => x"8c162283",
  5887 => x"dfff0655",
  5888 => x"748c1723",
  5889 => x"76800c89",
  5890 => x"3d0d04fa",
  5891 => x"3d0d788c",
  5892 => x"11227088",
  5893 => x"2a708106",
  5894 => x"51575856",
  5895 => x"74a9388c",
  5896 => x"162283df",
  5897 => x"ff065574",
  5898 => x"8c17237a",
  5899 => x"5479538e",
  5900 => x"16227090",
  5901 => x"2b70902c",
  5902 => x"545682c0",
  5903 => x"c0085256",
  5904 => x"83a73f88",
  5905 => x"3d0d0482",
  5906 => x"5480538e",
  5907 => x"16227090",
  5908 => x"2b70902c",
  5909 => x"545682c0",
  5910 => x"c0085257",
  5911 => x"85bd3f8c",
  5912 => x"162283df",
  5913 => x"ff065574",
  5914 => x"8c17237a",
  5915 => x"5479538e",
  5916 => x"16227090",
  5917 => x"2b70902c",
  5918 => x"545682c0",
  5919 => x"c0085256",
  5920 => x"82e73f88",
  5921 => x"3d0d04f9",
  5922 => x"3d0d797c",
  5923 => x"557b548e",
  5924 => x"11227090",
  5925 => x"2b70902c",
  5926 => x"555782c0",
  5927 => x"c0085358",
  5928 => x"5684f83f",
  5929 => x"80085780",
  5930 => x"08ff2e99",
  5931 => x"388c1622",
  5932 => x"a0800755",
  5933 => x"748c1723",
  5934 => x"800880d0",
  5935 => x"170c7680",
  5936 => x"0c893d0d",
  5937 => x"048c1622",
  5938 => x"83dfff06",
  5939 => x"55748c17",
  5940 => x"2376800c",
  5941 => x"893d0d04",
  5942 => x"fe3d0d74",
  5943 => x"8e112270",
  5944 => x"902b7090",
  5945 => x"2c555151",
  5946 => x"5382c0c0",
  5947 => x"085183c1",
  5948 => x"3f843d0d",
  5949 => x"04fb3d0d",
  5950 => x"77797072",
  5951 => x"07830653",
  5952 => x"54527093",
  5953 => x"38717373",
  5954 => x"08545654",
  5955 => x"7173082e",
  5956 => x"80c43873",
  5957 => x"75545271",
  5958 => x"337081ff",
  5959 => x"06525470",
  5960 => x"802e9d38",
  5961 => x"72335570",
  5962 => x"752e0981",
  5963 => x"06953881",
  5964 => x"12811471",
  5965 => x"337081ff",
  5966 => x"06545654",
  5967 => x"5270e538",
  5968 => x"72335573",
  5969 => x"81ff0675",
  5970 => x"81ff0671",
  5971 => x"7131800c",
  5972 => x"5252873d",
  5973 => x"0d047109",
  5974 => x"70f7fbfd",
  5975 => x"ff140670",
  5976 => x"f8848281",
  5977 => x"80065151",
  5978 => x"51709738",
  5979 => x"84148416",
  5980 => x"71085456",
  5981 => x"54717508",
  5982 => x"2edc3873",
  5983 => x"755452ff",
  5984 => x"9639800b",
  5985 => x"800c873d",
  5986 => x"0d04fd3d",
  5987 => x"0d757071",
  5988 => x"83065355",
  5989 => x"5270b838",
  5990 => x"71700870",
  5991 => x"09f7fbfd",
  5992 => x"ff120670",
  5993 => x"f8848281",
  5994 => x"80065151",
  5995 => x"5253709d",
  5996 => x"38841370",
  5997 => x"087009f7",
  5998 => x"fbfdff12",
  5999 => x"0670f884",
  6000 => x"82818006",
  6001 => x"51515253",
  6002 => x"70802ee5",
  6003 => x"38725271",
  6004 => x"33517080",
  6005 => x"2e8a3881",
  6006 => x"12703352",
  6007 => x"5270f838",
  6008 => x"71743180",
  6009 => x"0c853d0d",
  6010 => x"04fb3d0d",
  6011 => x"800b82d0",
  6012 => x"d40c7a53",
  6013 => x"79527851",
  6014 => x"84923f80",
  6015 => x"08558008",
  6016 => x"ff2e8838",
  6017 => x"74800c87",
  6018 => x"3d0d0482",
  6019 => x"d0d40856",
  6020 => x"75802ef0",
  6021 => x"38777671",
  6022 => x"0c547480",
  6023 => x"0c873d0d",
  6024 => x"04fb3d0d",
  6025 => x"787a2952",
  6026 => x"7751c9d9",
  6027 => x"3f800880",
  6028 => x"08555680",
  6029 => x"08802e80",
  6030 => x"e3388008",
  6031 => x"fc0508fc",
  6032 => x"06fc0555",
  6033 => x"74a42680",
  6034 => x"da389375",
  6035 => x"27bb3880",
  6036 => x"0b800870",
  6037 => x"8405800c",
  6038 => x"0c800854",
  6039 => x"80747084",
  6040 => x"05560c9b",
  6041 => x"7527a238",
  6042 => x"80747084",
  6043 => x"05560c80",
  6044 => x"74708405",
  6045 => x"560ca375",
  6046 => x"278f3880",
  6047 => x"74708405",
  6048 => x"560c8074",
  6049 => x"70840556",
  6050 => x"0c807470",
  6051 => x"8405560c",
  6052 => x"80747084",
  6053 => x"05560c80",
  6054 => x"740c7554",
  6055 => x"73800c87",
  6056 => x"3d0d0474",
  6057 => x"53805280",
  6058 => x"0851d7b1",
  6059 => x"3f7554ec",
  6060 => x"39fd3d0d",
  6061 => x"800b82d0",
  6062 => x"d40c7651",
  6063 => x"84d73f80",
  6064 => x"08538008",
  6065 => x"ff2e8838",
  6066 => x"72800c85",
  6067 => x"3d0d0482",
  6068 => x"d0d40854",
  6069 => x"73802ef0",
  6070 => x"38757471",
  6071 => x"0c527280",
  6072 => x"0c853d0d",
  6073 => x"04fc3d0d",
  6074 => x"800b82d0",
  6075 => x"d40c7852",
  6076 => x"775186bf",
  6077 => x"3f800854",
  6078 => x"8008ff2e",
  6079 => x"88387380",
  6080 => x"0c863d0d",
  6081 => x"0482d0d4",
  6082 => x"08557480",
  6083 => x"2ef03876",
  6084 => x"75710c53",
  6085 => x"73800c86",
  6086 => x"3d0d04fb",
  6087 => x"3d0d800b",
  6088 => x"82d0d40c",
  6089 => x"7a537952",
  6090 => x"7851849b",
  6091 => x"3f800855",
  6092 => x"8008ff2e",
  6093 => x"88387480",
  6094 => x"0c873d0d",
  6095 => x"0482d0d4",
  6096 => x"08567580",
  6097 => x"2ef03877",
  6098 => x"76710c54",
  6099 => x"74800c87",
  6100 => x"3d0d04fb",
  6101 => x"3d0d800b",
  6102 => x"82d0d40c",
  6103 => x"7a537952",
  6104 => x"785182a0",
  6105 => x"3f800855",
  6106 => x"8008ff2e",
  6107 => x"88387480",
  6108 => x"0c873d0d",
  6109 => x"0482d0d4",
  6110 => x"08567580",
  6111 => x"2ef03877",
  6112 => x"76710c54",
  6113 => x"74800c87",
  6114 => x"3d0d04fe",
  6115 => x"3d0d82d0",
  6116 => x"cc085170",
  6117 => x"8a3882d0",
  6118 => x"d87082d0",
  6119 => x"cc0c5170",
  6120 => x"75125252",
  6121 => x"ff537087",
  6122 => x"fb808026",
  6123 => x"88387082",
  6124 => x"d0cc0c71",
  6125 => x"5372800c",
  6126 => x"843d0d04",
  6127 => x"fd3d0d80",
  6128 => x"0b82c0b4",
  6129 => x"08545472",
  6130 => x"812e9e38",
  6131 => x"7382d0d0",
  6132 => x"0cfecad2",
  6133 => x"3ffec8a8",
  6134 => x"3f82d0a4",
  6135 => x"528151fe",
  6136 => x"c9e33f80",
  6137 => x"085185cb",
  6138 => x"3f7282d0",
  6139 => x"d00cfeca",
  6140 => x"b53ffec8",
  6141 => x"8b3f82d0",
  6142 => x"a4528151",
  6143 => x"fec9c63f",
  6144 => x"80085185",
  6145 => x"ae3f00ff",
  6146 => x"3900ff39",
  6147 => x"f53d0d7e",
  6148 => x"6082d0d0",
  6149 => x"08705b58",
  6150 => x"5b5b7580",
  6151 => x"c538777a",
  6152 => x"25a23877",
  6153 => x"1b703370",
  6154 => x"81ff0658",
  6155 => x"5859758a",
  6156 => x"2e993876",
  6157 => x"81ff0651",
  6158 => x"fec9cc3f",
  6159 => x"81185879",
  6160 => x"7824e038",
  6161 => x"79800c8d",
  6162 => x"3d0d048d",
  6163 => x"51fec9b7",
  6164 => x"3f783370",
  6165 => x"81ff0652",
  6166 => x"57fec9ab",
  6167 => x"3f811858",
  6168 => x"de397955",
  6169 => x"7a547d53",
  6170 => x"85528d3d",
  6171 => x"fc0551fe",
  6172 => x"c7d03f80",
  6173 => x"085684b4",
  6174 => x"3f7b8008",
  6175 => x"0c75800c",
  6176 => x"8d3d0d04",
  6177 => x"f63d0d7d",
  6178 => x"7f82d0d0",
  6179 => x"08705b58",
  6180 => x"5a5a7580",
  6181 => x"c4387779",
  6182 => x"25b638fe",
  6183 => x"c8c63f80",
  6184 => x"0881ff06",
  6185 => x"708d3270",
  6186 => x"30709f2a",
  6187 => x"51515757",
  6188 => x"768a2e80",
  6189 => x"c6387580",
  6190 => x"2e80c038",
  6191 => x"771a5676",
  6192 => x"76347651",
  6193 => x"fec8c03f",
  6194 => x"81185878",
  6195 => x"7824cc38",
  6196 => x"77567580",
  6197 => x"0c8c3d0d",
  6198 => x"04785579",
  6199 => x"547c5384",
  6200 => x"528c3dfc",
  6201 => x"0551fec6",
  6202 => x"d93f8008",
  6203 => x"5683bd3f",
  6204 => x"7a80080c",
  6205 => x"75800c8c",
  6206 => x"3d0d0477",
  6207 => x"1a568a76",
  6208 => x"34811858",
  6209 => x"8d51fec7",
  6210 => x"fe3f8a51",
  6211 => x"fec7f83f",
  6212 => x"7756ffbe",
  6213 => x"39fb3d0d",
  6214 => x"82d0d008",
  6215 => x"70565473",
  6216 => x"88387480",
  6217 => x"0c873d0d",
  6218 => x"04775383",
  6219 => x"52873dfc",
  6220 => x"0551fec6",
  6221 => x"8d3f8008",
  6222 => x"5482f13f",
  6223 => x"7580080c",
  6224 => x"73800c87",
  6225 => x"3d0d04fa",
  6226 => x"3d0d82d0",
  6227 => x"d008802e",
  6228 => x"a3387a55",
  6229 => x"79547853",
  6230 => x"8652883d",
  6231 => x"fc0551fe",
  6232 => x"c5e03f80",
  6233 => x"085682c4",
  6234 => x"3f768008",
  6235 => x"0c75800c",
  6236 => x"883d0d04",
  6237 => x"82b63f9d",
  6238 => x"0b80080c",
  6239 => x"ff0b800c",
  6240 => x"883d0d04",
  6241 => x"fb3d0d77",
  6242 => x"79565680",
  6243 => x"70545473",
  6244 => x"75259f38",
  6245 => x"74101010",
  6246 => x"f8055272",
  6247 => x"16703370",
  6248 => x"742b7607",
  6249 => x"8116f816",
  6250 => x"56565651",
  6251 => x"51747324",
  6252 => x"ea387380",
  6253 => x"0c873d0d",
  6254 => x"04fc3d0d",
  6255 => x"76785555",
  6256 => x"bc538052",
  6257 => x"7351d195",
  6258 => x"3f845274",
  6259 => x"51ffb53f",
  6260 => x"80087423",
  6261 => x"84528415",
  6262 => x"51ffa93f",
  6263 => x"80088215",
  6264 => x"23845288",
  6265 => x"1551ff9c",
  6266 => x"3f800884",
  6267 => x"150c8452",
  6268 => x"8c1551ff",
  6269 => x"8f3f8008",
  6270 => x"88152384",
  6271 => x"52901551",
  6272 => x"ff823f80",
  6273 => x"088a1523",
  6274 => x"84529415",
  6275 => x"51fef53f",
  6276 => x"80088c15",
  6277 => x"23845298",
  6278 => x"1551fee8",
  6279 => x"3f80088e",
  6280 => x"15238852",
  6281 => x"9c1551fe",
  6282 => x"db3f8008",
  6283 => x"90150c86",
  6284 => x"3d0d04e9",
  6285 => x"3d0d6a82",
  6286 => x"d0d00857",
  6287 => x"57759338",
  6288 => x"80c0800b",
  6289 => x"84180c75",
  6290 => x"ac180c75",
  6291 => x"800c993d",
  6292 => x"0d04893d",
  6293 => x"70556a54",
  6294 => x"558a5299",
  6295 => x"3dffbc05",
  6296 => x"51fec3de",
  6297 => x"3f800877",
  6298 => x"53755256",
  6299 => x"fecb3fbc",
  6300 => x"3f778008",
  6301 => x"0c75800c",
  6302 => x"993d0d04",
  6303 => x"fc3d0d81",
  6304 => x"5482d0d0",
  6305 => x"08883873",
  6306 => x"800c863d",
  6307 => x"0d047653",
  6308 => x"97b95286",
  6309 => x"3dfc0551",
  6310 => x"fec3a73f",
  6311 => x"8008548c",
  6312 => x"3f748008",
  6313 => x"0c73800c",
  6314 => x"863d0d04",
  6315 => x"82c0c008",
  6316 => x"800c04f7",
  6317 => x"3d0d7b82",
  6318 => x"c0c00882",
  6319 => x"c811085a",
  6320 => x"545a7780",
  6321 => x"2e80da38",
  6322 => x"81881884",
  6323 => x"1908ff05",
  6324 => x"81712b59",
  6325 => x"55598074",
  6326 => x"2480ea38",
  6327 => x"807424b5",
  6328 => x"3873822b",
  6329 => x"78118805",
  6330 => x"56568180",
  6331 => x"19087706",
  6332 => x"5372802e",
  6333 => x"b6387816",
  6334 => x"70085353",
  6335 => x"79517408",
  6336 => x"53722dff",
  6337 => x"14fc17fc",
  6338 => x"1779812c",
  6339 => x"5a575754",
  6340 => x"738025d6",
  6341 => x"38770858",
  6342 => x"77ffad38",
  6343 => x"82c0c008",
  6344 => x"53bc1308",
  6345 => x"a5387951",
  6346 => x"f9dc3f74",
  6347 => x"0853722d",
  6348 => x"ff14fc17",
  6349 => x"fc177981",
  6350 => x"2c5a5757",
  6351 => x"54738025",
  6352 => x"ffa838d1",
  6353 => x"398057ff",
  6354 => x"93397251",
  6355 => x"bc130853",
  6356 => x"722d7951",
  6357 => x"f9b03f8c",
  6358 => x"08028c0c",
  6359 => x"d43d0d8c",
  6360 => x"08880508",
  6361 => x"518e963f",
  6362 => x"80085473",
  6363 => x"802e9038",
  6364 => x"8c088805",
  6365 => x"08708c08",
  6366 => x"d0050c54",
  6367 => x"8cf5398c",
  6368 => x"088c0508",
  6369 => x"518df63f",
  6370 => x"80085473",
  6371 => x"802e9038",
  6372 => x"8c088c05",
  6373 => x"08708c08",
  6374 => x"d0050c54",
  6375 => x"8cd5398c",
  6376 => x"08880508",
  6377 => x"518da23f",
  6378 => x"80085473",
  6379 => x"802e80c5",
  6380 => x"388c088c",
  6381 => x"0508518d",
  6382 => x"903f8008",
  6383 => x"5473802e",
  6384 => x"a5388c08",
  6385 => x"8805088c",
  6386 => x"088c0508",
  6387 => x"55558415",
  6388 => x"08841508",
  6389 => x"2e90388c",
  6390 => x"db3f8008",
  6391 => x"708c08d0",
  6392 => x"050c548c",
  6393 => x"8e398c08",
  6394 => x"88050870",
  6395 => x"8c08d005",
  6396 => x"0c548bff",
  6397 => x"398c088c",
  6398 => x"0508518c",
  6399 => x"cc3f8008",
  6400 => x"5473802e",
  6401 => x"90388c08",
  6402 => x"8c050870",
  6403 => x"8c08d005",
  6404 => x"0c548bdf",
  6405 => x"398c088c",
  6406 => x"0508518b",
  6407 => x"e33f8008",
  6408 => x"5473802e",
  6409 => x"80e7388c",
  6410 => x"08880508",
  6411 => x"518bd13f",
  6412 => x"80085473",
  6413 => x"802e80c6",
  6414 => x"388c0890",
  6415 => x"05088c08",
  6416 => x"88050871",
  6417 => x"58565494",
  6418 => x"70547553",
  6419 => x"765254fe",
  6420 => x"c9bd3f8c",
  6421 => x"08900508",
  6422 => x"8c088805",
  6423 => x"088c088c",
  6424 => x"05088412",
  6425 => x"08841208",
  6426 => x"0684140c",
  6427 => x"8c089005",
  6428 => x"08708c08",
  6429 => x"d0050c51",
  6430 => x"5656568a",
  6431 => x"f6398c08",
  6432 => x"88050870",
  6433 => x"8c08d005",
  6434 => x"0c548ae7",
  6435 => x"398c0888",
  6436 => x"0508518a",
  6437 => x"eb3f8008",
  6438 => x"5473802e",
  6439 => x"90388c08",
  6440 => x"8c050870",
  6441 => x"8c08d005",
  6442 => x"0c548ac7",
  6443 => x"398c0888",
  6444 => x"05088811",
  6445 => x"088c08f4",
  6446 => x"050c8c08",
  6447 => x"8c050888",
  6448 => x"11088c08",
  6449 => x"f0050c8c",
  6450 => x"08880508",
  6451 => x"51515490",
  6452 => x"14088c15",
  6453 => x"08555573",
  6454 => x"8c08e805",
  6455 => x"0c748c08",
  6456 => x"ec050c8c",
  6457 => x"088c0508",
  6458 => x"54901408",
  6459 => x"8c150855",
  6460 => x"55738c08",
  6461 => x"e0050c74",
  6462 => x"8c08e405",
  6463 => x"0c8c08f4",
  6464 => x"05088c08",
  6465 => x"f0050831",
  6466 => x"8c08dc05",
  6467 => x"0c8c08dc",
  6468 => x"05088025",
  6469 => x"8c388c08",
  6470 => x"dc050830",
  6471 => x"8c08dc05",
  6472 => x"0c8c08dc",
  6473 => x"0508bf24",
  6474 => x"81b3388c",
  6475 => x"08f00508",
  6476 => x"8c08f405",
  6477 => x"082580cc",
  6478 => x"388c08f0",
  6479 => x"05088105",
  6480 => x"8c08f005",
  6481 => x"0c8c08e0",
  6482 => x"05088006",
  6483 => x"8c08e405",
  6484 => x"0881068c",
  6485 => x"08e00508",
  6486 => x"9f2b8c08",
  6487 => x"e4050881",
  6488 => x"2a707207",
  6489 => x"8c08e005",
  6490 => x"08812a70",
  6491 => x"76078c08",
  6492 => x"e0050c74",
  6493 => x"72078c08",
  6494 => x"e4050c59",
  6495 => x"595b5b58",
  6496 => x"56ffa839",
  6497 => x"8c08f405",
  6498 => x"088c08f0",
  6499 => x"05082581",
  6500 => x"8f388c08",
  6501 => x"f4050881",
  6502 => x"058c08f4",
  6503 => x"050c8c08",
  6504 => x"e8050880",
  6505 => x"068c08ec",
  6506 => x"05088106",
  6507 => x"8c08e805",
  6508 => x"089f2b8c",
  6509 => x"08ec0508",
  6510 => x"812a7072",
  6511 => x"078c08e8",
  6512 => x"0508812a",
  6513 => x"7076078c",
  6514 => x"08e8050c",
  6515 => x"7472078c",
  6516 => x"08ec050c",
  6517 => x"59595b5b",
  6518 => x"5856ffa8",
  6519 => x"398c08f0",
  6520 => x"05088c08",
  6521 => x"f4050825",
  6522 => x"9d388c08",
  6523 => x"f405088c",
  6524 => x"08f0050c",
  6525 => x"80548055",
  6526 => x"738c08e0",
  6527 => x"050c748c",
  6528 => x"08e4050c",
  6529 => x"9b398c08",
  6530 => x"f005088c",
  6531 => x"08f4050c",
  6532 => x"80548055",
  6533 => x"738c08e8",
  6534 => x"050c748c",
  6535 => x"08ec050c",
  6536 => x"8c088805",
  6537 => x"088c088c",
  6538 => x"05085555",
  6539 => x"84150884",
  6540 => x"15082e84",
  6541 => x"e5388c08",
  6542 => x"88050854",
  6543 => x"84140880",
  6544 => x"2e81b538",
  6545 => x"8c08e005",
  6546 => x"088c08e4",
  6547 => x"05085654",
  6548 => x"738c08c8",
  6549 => x"050c748c",
  6550 => x"08cc050c",
  6551 => x"8c08e805",
  6552 => x"088c08ec",
  6553 => x"05085755",
  6554 => x"748c08c0",
  6555 => x"050c758c",
  6556 => x"08c4050c",
  6557 => x"8c08cc05",
  6558 => x"088c08c4",
  6559 => x"05087171",
  6560 => x"31708c08",
  6561 => x"ffbc050c",
  6562 => x"52555681",
  6563 => x"0b8c08ff",
  6564 => x"b4050c8c",
  6565 => x"08ffbc05",
  6566 => x"088c08cc",
  6567 => x"05085755",
  6568 => x"74762689",
  6569 => x"38800b8c",
  6570 => x"08ffb405",
  6571 => x"0c8c08c8",
  6572 => x"05088c08",
  6573 => x"c0050871",
  6574 => x"7131708c",
  6575 => x"08ffb805",
  6576 => x"0c8c08ff",
  6577 => x"b8050870",
  6578 => x"8c08ffb4",
  6579 => x"05083170",
  6580 => x"8c08ffb8",
  6581 => x"050c5259",
  6582 => x"5256548c",
  6583 => x"08ffb805",
  6584 => x"088c08ff",
  6585 => x"bc050856",
  6586 => x"54738c08",
  6587 => x"f8050c74",
  6588 => x"8c08fc05",
  6589 => x"0c81bb39",
  6590 => x"8c08e805",
  6591 => x"088c08ec",
  6592 => x"05085755",
  6593 => x"748c08ff",
  6594 => x"ac050c75",
  6595 => x"8c08ffb0",
  6596 => x"050c8c08",
  6597 => x"e005088c",
  6598 => x"08e40508",
  6599 => x"5654738c",
  6600 => x"08ffa405",
  6601 => x"0c748c08",
  6602 => x"ffa8050c",
  6603 => x"8c08ffb0",
  6604 => x"05088c08",
  6605 => x"ffa80508",
  6606 => x"71713170",
  6607 => x"8c08ffa0",
  6608 => x"050c5257",
  6609 => x"55810b8c",
  6610 => x"08ff9805",
  6611 => x"0c8c08ff",
  6612 => x"a005088c",
  6613 => x"08ffb005",
  6614 => x"08565473",
  6615 => x"75268938",
  6616 => x"800b8c08",
  6617 => x"ff98050c",
  6618 => x"8c08ffac",
  6619 => x"05088c08",
  6620 => x"ffa40508",
  6621 => x"71713170",
  6622 => x"8c08ff9c",
  6623 => x"050c8c08",
  6624 => x"ff9c0508",
  6625 => x"708c08ff",
  6626 => x"98050831",
  6627 => x"708c08ff",
  6628 => x"9c050c53",
  6629 => x"58525556",
  6630 => x"8c08ff9c",
  6631 => x"05088c08",
  6632 => x"ffa00508",
  6633 => x"5654738c",
  6634 => x"08f8050c",
  6635 => x"748c08fc",
  6636 => x"050c800b",
  6637 => x"8c08f805",
  6638 => x"0824b738",
  6639 => x"8c089005",
  6640 => x"0854800b",
  6641 => x"84150c8c",
  6642 => x"08900508",
  6643 => x"8c08f405",
  6644 => x"0888120c",
  6645 => x"8c089005",
  6646 => x"0857548c",
  6647 => x"08f80508",
  6648 => x"8c08fc05",
  6649 => x"08565473",
  6650 => x"8c170c74",
  6651 => x"90170c80",
  6652 => x"cf398c08",
  6653 => x"90050854",
  6654 => x"810b8415",
  6655 => x"0c8c0890",
  6656 => x"05088c08",
  6657 => x"f4050888",
  6658 => x"120c8c08",
  6659 => x"9005088c",
  6660 => x"08d40558",
  6661 => x"58548c08",
  6662 => x"f805088c",
  6663 => x"08fc0508",
  6664 => x"56547352",
  6665 => x"74537551",
  6666 => x"80c8c93f",
  6667 => x"8c08d405",
  6668 => x"088c08d8",
  6669 => x"05085654",
  6670 => x"738c180c",
  6671 => x"7490180c",
  6672 => x"8c089005",
  6673 => x"08548c14",
  6674 => x"08f00a26",
  6675 => x"82b1388c",
  6676 => x"08900508",
  6677 => x"8c110870",
  6678 => x"90130807",
  6679 => x"51555573",
  6680 => x"802e829b",
  6681 => x"388c0890",
  6682 => x"05088c08",
  6683 => x"90050890",
  6684 => x"11089f2a",
  6685 => x"8c120810",
  6686 => x"7072078c",
  6687 => x"150c9013",
  6688 => x"08109015",
  6689 => x"0c8c0890",
  6690 => x"05088811",
  6691 => x"08ff0588",
  6692 => x"120c5358",
  6693 => x"585557ff",
  6694 => x"a7398c08",
  6695 => x"9005088c",
  6696 => x"08880508",
  6697 => x"84110884",
  6698 => x"130c8c08",
  6699 => x"9005088c",
  6700 => x"08f40508",
  6701 => x"88120c8c",
  6702 => x"08900508",
  6703 => x"8c08ff94",
  6704 => x"050c5256",
  6705 => x"548c08e8",
  6706 => x"05088c08",
  6707 => x"ec050857",
  6708 => x"55748c08",
  6709 => x"ff8c050c",
  6710 => x"758c08ff",
  6711 => x"90050c8c",
  6712 => x"08e00508",
  6713 => x"8c08e405",
  6714 => x"08565473",
  6715 => x"8c08ff84",
  6716 => x"050c748c",
  6717 => x"08ff8805",
  6718 => x"0c8c08ff",
  6719 => x"9005088c",
  6720 => x"08ff8805",
  6721 => x"08701270",
  6722 => x"8c08ff80",
  6723 => x"050c5257",
  6724 => x"55810b8c",
  6725 => x"08fef805",
  6726 => x"0c8c08ff",
  6727 => x"8005088c",
  6728 => x"08ff9005",
  6729 => x"08565474",
  6730 => x"74268938",
  6731 => x"800b8c08",
  6732 => x"fef8050c",
  6733 => x"8c08ff8c",
  6734 => x"05088c08",
  6735 => x"ff840508",
  6736 => x"7012708c",
  6737 => x"08fefc05",
  6738 => x"0c8c08fe",
  6739 => x"fc05088c",
  6740 => x"08fef805",
  6741 => x"0811708c",
  6742 => x"08fefc05",
  6743 => x"0c535852",
  6744 => x"55568c08",
  6745 => x"fefc0508",
  6746 => x"8c08ff80",
  6747 => x"05088c08",
  6748 => x"ff940508",
  6749 => x"58565473",
  6750 => x"8c170c74",
  6751 => x"90170c8c",
  6752 => x"08900508",
  6753 => x"5483740c",
  6754 => x"8c089005",
  6755 => x"08548c14",
  6756 => x"08f80a26",
  6757 => x"843880cf",
  6758 => x"398c0890",
  6759 => x"05088c08",
  6760 => x"9005088c",
  6761 => x"11088006",
  6762 => x"90120881",
  6763 => x"068c0890",
  6764 => x"05088c11",
  6765 => x"089f2b90",
  6766 => x"1208812a",
  6767 => x"7072078c",
  6768 => x"1408812a",
  6769 => x"7077078c",
  6770 => x"1a0c7572",
  6771 => x"07901a0c",
  6772 => x"8c089005",
  6773 => x"08881108",
  6774 => x"81058812",
  6775 => x"0c51575c",
  6776 => x"5f5f5c5a",
  6777 => x"58555b8c",
  6778 => x"08900508",
  6779 => x"708c08d0",
  6780 => x"050c548c",
  6781 => x"08d00508",
  6782 => x"800cae3d",
  6783 => x"0d8c0c04",
  6784 => x"8c08028c",
  6785 => x"0cff3d0d",
  6786 => x"800b8c08",
  6787 => x"fc050c8c",
  6788 => x"08880508",
  6789 => x"51700882",
  6790 => x"2e098106",
  6791 => x"8838810b",
  6792 => x"8c08fc05",
  6793 => x"0c8c08fc",
  6794 => x"05087080",
  6795 => x"0c51833d",
  6796 => x"0d8c0c04",
  6797 => x"8c08028c",
  6798 => x"0c803d0d",
  6799 => x"82c08c70",
  6800 => x"800c5182",
  6801 => x"3d0d8c0c",
  6802 => x"048c0802",
  6803 => x"8c0cff3d",
  6804 => x"0d800b8c",
  6805 => x"08fc050c",
  6806 => x"8c088805",
  6807 => x"08517008",
  6808 => x"842e0981",
  6809 => x"06883881",
  6810 => x"0b8c08fc",
  6811 => x"050c8c08",
  6812 => x"fc050870",
  6813 => x"800c5183",
  6814 => x"3d0d8c0c",
  6815 => x"048c0802",
  6816 => x"8c0cff3d",
  6817 => x"0d800b8c",
  6818 => x"08fc050c",
  6819 => x"8c088805",
  6820 => x"08517008",
  6821 => x"802e8f38",
  6822 => x"8c088805",
  6823 => x"08517008",
  6824 => x"812e8338",
  6825 => x"8839810b",
  6826 => x"8c08fc05",
  6827 => x"0c8c08fc",
  6828 => x"05087080",
  6829 => x"0c51833d",
  6830 => x"0d8c0c04",
  6831 => x"8c08028c",
  6832 => x"0ce73d0d",
  6833 => x"8c088805",
  6834 => x"08568c08",
  6835 => x"8c05088c",
  6836 => x"08900508",
  6837 => x"5654738c",
  6838 => x"08ffb805",
  6839 => x"0c748c08",
  6840 => x"ffbc050c",
  6841 => x"8c089405",
  6842 => x"088c0898",
  6843 => x"05085654",
  6844 => x"738c08ff",
  6845 => x"b0050c74",
  6846 => x"8c08ffb4",
  6847 => x"050c8c08",
  6848 => x"ec057053",
  6849 => x"8c08ffb8",
  6850 => x"05705351",
  6851 => x"5480d6be",
  6852 => x"3f8c08d8",
  6853 => x"0570538c",
  6854 => x"08ffb005",
  6855 => x"70535154",
  6856 => x"80d6ab3f",
  6857 => x"8c08c405",
  6858 => x"70548c08",
  6859 => x"d8057054",
  6860 => x"8c08ec05",
  6861 => x"70545151",
  6862 => x"54f09c3f",
  6863 => x"8008708c",
  6864 => x"08c0050c",
  6865 => x"8c08c005",
  6866 => x"08537652",
  6867 => x"5480c5c8",
  6868 => x"3f75800c",
  6869 => x"9b3d0d8c",
  6870 => x"0c048c08",
  6871 => x"028c0ce7",
  6872 => x"3d0d8c08",
  6873 => x"88050856",
  6874 => x"8c088c05",
  6875 => x"088c0890",
  6876 => x"05085654",
  6877 => x"738c08ff",
  6878 => x"b8050c74",
  6879 => x"8c08ffbc",
  6880 => x"050c8c08",
  6881 => x"9405088c",
  6882 => x"08980508",
  6883 => x"5654738c",
  6884 => x"08ffb005",
  6885 => x"0c748c08",
  6886 => x"ffb4050c",
  6887 => x"8c08ec05",
  6888 => x"70538c08",
  6889 => x"ffb80570",
  6890 => x"53515480",
  6891 => x"d5a03f8c",
  6892 => x"08d80570",
  6893 => x"538c08ff",
  6894 => x"b0057053",
  6895 => x"515480d5",
  6896 => x"8d3f8c08",
  6897 => x"dc050881",
  6898 => x"328c08dc",
  6899 => x"050c8c08",
  6900 => x"c4057054",
  6901 => x"8c08d805",
  6902 => x"70548c08",
  6903 => x"ec057054",
  6904 => x"515154ee",
  6905 => x"f23f8008",
  6906 => x"708c08c0",
  6907 => x"050c8c08",
  6908 => x"c0050853",
  6909 => x"76525480",
  6910 => x"c49e3f75",
  6911 => x"800c9b3d",
  6912 => x"0d8c0c04",
  6913 => x"8c08028c",
  6914 => x"0cff833d",
  6915 => x"0d8c088c",
  6916 => x"05088c08",
  6917 => x"90050858",
  6918 => x"56758c08",
  6919 => x"ffb8050c",
  6920 => x"768c08ff",
  6921 => x"bc050c8c",
  6922 => x"08940508",
  6923 => x"8c089805",
  6924 => x"08585675",
  6925 => x"8c08ffb0",
  6926 => x"050c768c",
  6927 => x"08ffb405",
  6928 => x"0c8c08ec",
  6929 => x"0570538c",
  6930 => x"08ffb805",
  6931 => x"70535156",
  6932 => x"80d3fb3f",
  6933 => x"8c08d805",
  6934 => x"70538c08",
  6935 => x"ffb00570",
  6936 => x"53515680",
  6937 => x"d3e83f8c",
  6938 => x"08ec058c",
  6939 => x"08ffac05",
  6940 => x"0c8c08d8",
  6941 => x"058c08ff",
  6942 => x"a8050c8c",
  6943 => x"08c4058c",
  6944 => x"08ffa405",
  6945 => x"0c805680",
  6946 => x"57758c08",
  6947 => x"ff98050c",
  6948 => x"768c08ff",
  6949 => x"9c050c80",
  6950 => x"56805775",
  6951 => x"8c08ff90",
  6952 => x"050c768c",
  6953 => x"08ff9405",
  6954 => x"0c8c08ff",
  6955 => x"ac050851",
  6956 => x"9ba23f80",
  6957 => x"08567580",
  6958 => x"2e80d338",
  6959 => x"8c08ffac",
  6960 => x"05088c08",
  6961 => x"fec4050c",
  6962 => x"800b8c08",
  6963 => x"fec0050c",
  6964 => x"8c08ffac",
  6965 => x"05088c08",
  6966 => x"ffa80508",
  6967 => x"57578417",
  6968 => x"08841708",
  6969 => x"2e893881",
  6970 => x"0b8c08fe",
  6971 => x"c0050c8c",
  6972 => x"08fec405",
  6973 => x"088c08fe",
  6974 => x"c0050884",
  6975 => x"120c8c08",
  6976 => x"ffac0508",
  6977 => x"8c08ffa0",
  6978 => x"050c5699",
  6979 => x"a0398c08",
  6980 => x"ffa80508",
  6981 => x"519abd3f",
  6982 => x"80085675",
  6983 => x"802e80d3",
  6984 => x"388c08ff",
  6985 => x"a805088c",
  6986 => x"08febc05",
  6987 => x"0c800b8c",
  6988 => x"08feb805",
  6989 => x"0c8c08ff",
  6990 => x"ac05088c",
  6991 => x"08ffa805",
  6992 => x"08575784",
  6993 => x"17088417",
  6994 => x"082e8938",
  6995 => x"810b8c08",
  6996 => x"feb8050c",
  6997 => x"8c08febc",
  6998 => x"05088c08",
  6999 => x"feb80508",
  7000 => x"84120c8c",
  7001 => x"08ffa805",
  7002 => x"088c08ff",
  7003 => x"a0050c57",
  7004 => x"98bb398c",
  7005 => x"08ffac05",
  7006 => x"085199a4",
  7007 => x"3f800856",
  7008 => x"75802e80",
  7009 => x"f5388c08",
  7010 => x"ffa80508",
  7011 => x"5198dd3f",
  7012 => x"80085675",
  7013 => x"802e9138",
  7014 => x"98bd3f80",
  7015 => x"08708c08",
  7016 => x"ffa0050c",
  7017 => x"56988639",
  7018 => x"8c08ffac",
  7019 => x"05088c08",
  7020 => x"feb4050c",
  7021 => x"800b8c08",
  7022 => x"feb0050c",
  7023 => x"8c08ffac",
  7024 => x"05088c08",
  7025 => x"ffa80508",
  7026 => x"57578417",
  7027 => x"08841708",
  7028 => x"2e893881",
  7029 => x"0b8c08fe",
  7030 => x"b0050c8c",
  7031 => x"08feb405",
  7032 => x"088c08fe",
  7033 => x"b0050884",
  7034 => x"120c8c08",
  7035 => x"ffac0508",
  7036 => x"8c08ffa0",
  7037 => x"050c5697",
  7038 => x"b4398c08",
  7039 => x"ffa80508",
  7040 => x"51989d3f",
  7041 => x"80085675",
  7042 => x"802e80f5",
  7043 => x"388c08ff",
  7044 => x"ac050851",
  7045 => x"97d63f80",
  7046 => x"08567580",
  7047 => x"2e913897",
  7048 => x"b63f8008",
  7049 => x"708c08ff",
  7050 => x"a0050c56",
  7051 => x"96ff398c",
  7052 => x"08ffa805",
  7053 => x"088c08fe",
  7054 => x"ac050c80",
  7055 => x"0b8c08fe",
  7056 => x"a8050c8c",
  7057 => x"08ffac05",
  7058 => x"088c08ff",
  7059 => x"a8050857",
  7060 => x"57841708",
  7061 => x"8417082e",
  7062 => x"8938810b",
  7063 => x"8c08fea8",
  7064 => x"050c8c08",
  7065 => x"feac0508",
  7066 => x"8c08fea8",
  7067 => x"05088412",
  7068 => x"0c8c08ff",
  7069 => x"a805088c",
  7070 => x"08ffa005",
  7071 => x"0c5796ad",
  7072 => x"398c08ff",
  7073 => x"ac050851",
  7074 => x"96e23f80",
  7075 => x"08567580",
  7076 => x"2e80d338",
  7077 => x"8c08ffac",
  7078 => x"05088c08",
  7079 => x"fea4050c",
  7080 => x"800b8c08",
  7081 => x"fea0050c",
  7082 => x"8c08ffac",
  7083 => x"05088c08",
  7084 => x"ffa80508",
  7085 => x"57578417",
  7086 => x"08841708",
  7087 => x"2e893881",
  7088 => x"0b8c08fe",
  7089 => x"a0050c8c",
  7090 => x"08fea405",
  7091 => x"088c08fe",
  7092 => x"a0050884",
  7093 => x"120c8c08",
  7094 => x"ffac0508",
  7095 => x"8c08ffa0",
  7096 => x"050c5695",
  7097 => x"c8398c08",
  7098 => x"ffa80508",
  7099 => x"5195fd3f",
  7100 => x"80085675",
  7101 => x"802e80d3",
  7102 => x"388c08ff",
  7103 => x"a805088c",
  7104 => x"08fe9c05",
  7105 => x"0c800b8c",
  7106 => x"08fe9805",
  7107 => x"0c8c08ff",
  7108 => x"ac05088c",
  7109 => x"08ffa805",
  7110 => x"08575784",
  7111 => x"17088417",
  7112 => x"082e8938",
  7113 => x"810b8c08",
  7114 => x"fe98050c",
  7115 => x"8c08fe9c",
  7116 => x"05088c08",
  7117 => x"fe980508",
  7118 => x"84120c8c",
  7119 => x"08ffa805",
  7120 => x"088c08ff",
  7121 => x"a0050c57",
  7122 => x"94e3398c",
  7123 => x"08ffac05",
  7124 => x"08901108",
  7125 => x"8c08ff8c",
  7126 => x"050c8c08",
  7127 => x"ffac0508",
  7128 => x"8c110880",
  7129 => x"2a595956",
  7130 => x"80778c08",
  7131 => x"ff88050c",
  7132 => x"8c08ffa8",
  7133 => x"05089011",
  7134 => x"088c08ff",
  7135 => x"84050c8c",
  7136 => x"08ffa805",
  7137 => x"088c1108",
  7138 => x"802a5a5a",
  7139 => x"51568077",
  7140 => x"8c08ff80",
  7141 => x"050c8c08",
  7142 => x"ff840508",
  7143 => x"5a56800b",
  7144 => x"8c08ff8c",
  7145 => x"05085858",
  7146 => x"800b8c08",
  7147 => x"fef0055b",
  7148 => x"56755476",
  7149 => x"55775278",
  7150 => x"537951b5",
  7151 => x"d93f8c08",
  7152 => x"fef00508",
  7153 => x"8c08fef4",
  7154 => x"05085856",
  7155 => x"758c08fe",
  7156 => x"f8050c76",
  7157 => x"8c08fefc",
  7158 => x"050c8c08",
  7159 => x"ff800508",
  7160 => x"59800b8c",
  7161 => x"08ff8c05",
  7162 => x"08585880",
  7163 => x"0b8c08fe",
  7164 => x"e8055b56",
  7165 => x"75547655",
  7166 => x"77527853",
  7167 => x"7951b596",
  7168 => x"3f8c08fe",
  7169 => x"e805088c",
  7170 => x"08feec05",
  7171 => x"08585675",
  7172 => x"8c08fef0",
  7173 => x"050c768c",
  7174 => x"08fef405",
  7175 => x"0c8c08ff",
  7176 => x"84050859",
  7177 => x"800b8c08",
  7178 => x"ff880508",
  7179 => x"5858800b",
  7180 => x"8c08fee0",
  7181 => x"055b5675",
  7182 => x"54765577",
  7183 => x"52785379",
  7184 => x"51b4d33f",
  7185 => x"8c08fee0",
  7186 => x"05088c08",
  7187 => x"fee40508",
  7188 => x"5856758c",
  7189 => x"08fee805",
  7190 => x"0c768c08",
  7191 => x"feec050c",
  7192 => x"8c08ff80",
  7193 => x"05085980",
  7194 => x"0b8c08ff",
  7195 => x"88050858",
  7196 => x"58800b8c",
  7197 => x"08fed805",
  7198 => x"5b567554",
  7199 => x"76557752",
  7200 => x"78537951",
  7201 => x"b4903f8c",
  7202 => x"08fed805",
  7203 => x"088c08fe",
  7204 => x"dc050858",
  7205 => x"56758c08",
  7206 => x"fee0050c",
  7207 => x"768c08fe",
  7208 => x"e4050c80",
  7209 => x"56805775",
  7210 => x"8c08fed8",
  7211 => x"050c768c",
  7212 => x"08fedc05",
  7213 => x"0c805680",
  7214 => x"57758c08",
  7215 => x"fed0050c",
  7216 => x"768c08fe",
  7217 => x"d4050c8c",
  7218 => x"08fef005",
  7219 => x"088c08fe",
  7220 => x"f4050858",
  7221 => x"56758c08",
  7222 => x"fe90050c",
  7223 => x"768c08fe",
  7224 => x"94050c8c",
  7225 => x"08fee805",
  7226 => x"088c08fe",
  7227 => x"ec050858",
  7228 => x"56758c08",
  7229 => x"fe88050c",
  7230 => x"768c08fe",
  7231 => x"8c050c8c",
  7232 => x"08fe9405",
  7233 => x"088c08fe",
  7234 => x"8c050870",
  7235 => x"12708c08",
  7236 => x"fe84050c",
  7237 => x"52575781",
  7238 => x"0b8c08fd",
  7239 => x"fc050c8c",
  7240 => x"08fe8405",
  7241 => x"088c08fe",
  7242 => x"94050857",
  7243 => x"57757726",
  7244 => x"8938800b",
  7245 => x"8c08fdfc",
  7246 => x"050c8c08",
  7247 => x"fe900508",
  7248 => x"8c08fe88",
  7249 => x"05087012",
  7250 => x"708c08fe",
  7251 => x"80050c8c",
  7252 => x"08fe8005",
  7253 => x"088c08fd",
  7254 => x"fc050811",
  7255 => x"708c08fe",
  7256 => x"80050c53",
  7257 => x"51525757",
  7258 => x"8c08fe80",
  7259 => x"05088c08",
  7260 => x"fe840508",
  7261 => x"5856758c",
  7262 => x"08fec805",
  7263 => x"0c768c08",
  7264 => x"fecc050c",
  7265 => x"8c08fef0",
  7266 => x"05088c08",
  7267 => x"fec80508",
  7268 => x"26a6388c",
  7269 => x"08fef005",
  7270 => x"088c08fe",
  7271 => x"c805082e",
  7272 => x"09810681",
  7273 => x"c6388c08",
  7274 => x"fef40508",
  7275 => x"8c08fecc",
  7276 => x"05082684",
  7277 => x"3881b439",
  7278 => x"8c08fed8",
  7279 => x"05088c08",
  7280 => x"fedc0508",
  7281 => x"5856758c",
  7282 => x"08fdf405",
  7283 => x"0c768c08",
  7284 => x"fdf8050c",
  7285 => x"81568057",
  7286 => x"758c08fd",
  7287 => x"ec050c76",
  7288 => x"8c08fdf0",
  7289 => x"050c8c08",
  7290 => x"fdf80508",
  7291 => x"8c08fdf0",
  7292 => x"05087012",
  7293 => x"708c08fd",
  7294 => x"e8050c52",
  7295 => x"5757810b",
  7296 => x"8c08fde0",
  7297 => x"050c8c08",
  7298 => x"fde80508",
  7299 => x"8c08fdf8",
  7300 => x"05085757",
  7301 => x"75772689",
  7302 => x"38800b8c",
  7303 => x"08fde005",
  7304 => x"0c8c08fd",
  7305 => x"f405088c",
  7306 => x"08fdec05",
  7307 => x"08701270",
  7308 => x"8c08fde4",
  7309 => x"050c8c08",
  7310 => x"fde40508",
  7311 => x"8c08fde0",
  7312 => x"05081170",
  7313 => x"8c08fde4",
  7314 => x"050c5351",
  7315 => x"5257578c",
  7316 => x"08fde405",
  7317 => x"088c08fd",
  7318 => x"e8050858",
  7319 => x"56758c08",
  7320 => x"fed8050c",
  7321 => x"768c08fe",
  7322 => x"dc050c8c",
  7323 => x"08fecc05",
  7324 => x"08578077",
  7325 => x"802b8c08",
  7326 => x"fef0050c",
  7327 => x"56800b8c",
  7328 => x"08fef405",
  7329 => x"0c8c08fe",
  7330 => x"f805088c",
  7331 => x"08fefc05",
  7332 => x"08585675",
  7333 => x"8c08fdd8",
  7334 => x"050c768c",
  7335 => x"08fddc05",
  7336 => x"0c8c08fe",
  7337 => x"f005088c",
  7338 => x"08fef405",
  7339 => x"08585675",
  7340 => x"8c08fdd0",
  7341 => x"050c768c",
  7342 => x"08fdd405",
  7343 => x"0c8c08fd",
  7344 => x"dc05088c",
  7345 => x"08fdd405",
  7346 => x"08701270",
  7347 => x"8c08fdcc",
  7348 => x"050c5257",
  7349 => x"57810b8c",
  7350 => x"08fdc405",
  7351 => x"0c8c08fd",
  7352 => x"cc05088c",
  7353 => x"08fddc05",
  7354 => x"08575775",
  7355 => x"77268938",
  7356 => x"800b8c08",
  7357 => x"fdc4050c",
  7358 => x"8c08fdd8",
  7359 => x"05088c08",
  7360 => x"fdd00508",
  7361 => x"7012708c",
  7362 => x"08fdc805",
  7363 => x"0c8c08fd",
  7364 => x"c805088c",
  7365 => x"08fdc405",
  7366 => x"0811708c",
  7367 => x"08fdc805",
  7368 => x"0c535152",
  7369 => x"57578c08",
  7370 => x"fdc80508",
  7371 => x"8c08fdcc",
  7372 => x"05085856",
  7373 => x"758c08fe",
  7374 => x"d0050c76",
  7375 => x"8c08fed4",
  7376 => x"050c8c08",
  7377 => x"fef80508",
  7378 => x"8c08fed0",
  7379 => x"050826a6",
  7380 => x"388c08fe",
  7381 => x"f805088c",
  7382 => x"08fed005",
  7383 => x"082e0981",
  7384 => x"0681c638",
  7385 => x"8c08fefc",
  7386 => x"05088c08",
  7387 => x"fed40508",
  7388 => x"26843881",
  7389 => x"b4398c08",
  7390 => x"fed80508",
  7391 => x"8c08fedc",
  7392 => x"05085856",
  7393 => x"758c08fd",
  7394 => x"bc050c76",
  7395 => x"8c08fdc0",
  7396 => x"050c8056",
  7397 => x"8157758c",
  7398 => x"08fdb405",
  7399 => x"0c768c08",
  7400 => x"fdb8050c",
  7401 => x"8c08fdc0",
  7402 => x"05088c08",
  7403 => x"fdb80508",
  7404 => x"7012708c",
  7405 => x"08fdb005",
  7406 => x"0c525757",
  7407 => x"810b8c08",
  7408 => x"fda8050c",
  7409 => x"8c08fdb0",
  7410 => x"05088c08",
  7411 => x"fdc00508",
  7412 => x"57577577",
  7413 => x"26893880",
  7414 => x"0b8c08fd",
  7415 => x"a8050c8c",
  7416 => x"08fdbc05",
  7417 => x"088c08fd",
  7418 => x"b4050870",
  7419 => x"12708c08",
  7420 => x"fdac050c",
  7421 => x"8c08fdac",
  7422 => x"05088c08",
  7423 => x"fda80508",
  7424 => x"11708c08",
  7425 => x"fdac050c",
  7426 => x"53515257",
  7427 => x"578c08fd",
  7428 => x"ac05088c",
  7429 => x"08fdb005",
  7430 => x"08585675",
  7431 => x"8c08fed8",
  7432 => x"050c768c",
  7433 => x"08fedc05",
  7434 => x"0c8c08fe",
  7435 => x"c8050880",
  7436 => x"2a708c08",
  7437 => x"fda4050c",
  7438 => x"5780708c",
  7439 => x"08fda005",
  7440 => x"0c568c08",
  7441 => x"fda00508",
  7442 => x"8c08fda4",
  7443 => x"05085856",
  7444 => x"758c08fd",
  7445 => x"a0050c76",
  7446 => x"8c08fda4",
  7447 => x"050c8c08",
  7448 => x"fee00508",
  7449 => x"8c08fee4",
  7450 => x"05085856",
  7451 => x"758c08fd",
  7452 => x"98050c76",
  7453 => x"8c08fd9c",
  7454 => x"050c8c08",
  7455 => x"fda40508",
  7456 => x"8c08fd9c",
  7457 => x"05087012",
  7458 => x"708c08fd",
  7459 => x"94050c52",
  7460 => x"5757810b",
  7461 => x"8c08fd8c",
  7462 => x"050c8c08",
  7463 => x"fd940508",
  7464 => x"8c08fda4",
  7465 => x"05085757",
  7466 => x"75772689",
  7467 => x"38800b8c",
  7468 => x"08fd8c05",
  7469 => x"0c8c08fd",
  7470 => x"a005088c",
  7471 => x"08fd9805",
  7472 => x"08701270",
  7473 => x"8c08fd90",
  7474 => x"050c8c08",
  7475 => x"fd900508",
  7476 => x"8c08fd8c",
  7477 => x"05081170",
  7478 => x"8c08fd90",
  7479 => x"050c5351",
  7480 => x"5257578c",
  7481 => x"08fed805",
  7482 => x"088c08fe",
  7483 => x"dc050858",
  7484 => x"56758c08",
  7485 => x"fd84050c",
  7486 => x"768c08fd",
  7487 => x"88050c8c",
  7488 => x"08fd8805",
  7489 => x"088c08fd",
  7490 => x"94050870",
  7491 => x"12708c08",
  7492 => x"fd80050c",
  7493 => x"52575781",
  7494 => x"0b8c08fc",
  7495 => x"f8050c8c",
  7496 => x"08fd8005",
  7497 => x"088c08fd",
  7498 => x"88050857",
  7499 => x"57757726",
  7500 => x"8938800b",
  7501 => x"8c08fcf8",
  7502 => x"050c8c08",
  7503 => x"fd840508",
  7504 => x"8c08fd90",
  7505 => x"05087012",
  7506 => x"708c08fc",
  7507 => x"fc050c8c",
  7508 => x"08fcfc05",
  7509 => x"088c08fc",
  7510 => x"f8050811",
  7511 => x"708c08fc",
  7512 => x"fc050c53",
  7513 => x"51525757",
  7514 => x"8c08fcfc",
  7515 => x"05088c08",
  7516 => x"fd800508",
  7517 => x"5856758c",
  7518 => x"08fed805",
  7519 => x"0c768c08",
  7520 => x"fedc050c",
  7521 => x"8c08fed8",
  7522 => x"05088c08",
  7523 => x"fedc0508",
  7524 => x"5856758c",
  7525 => x"08ff9005",
  7526 => x"0c768c08",
  7527 => x"ff94050c",
  7528 => x"8c08fed0",
  7529 => x"05088c08",
  7530 => x"fed40508",
  7531 => x"5856758c",
  7532 => x"08ff9805",
  7533 => x"0c768c08",
  7534 => x"ff9c050c",
  7535 => x"8c08ffa4",
  7536 => x"05088c08",
  7537 => x"ffac0508",
  7538 => x"8c08ffa8",
  7539 => x"05088812",
  7540 => x"08881208",
  7541 => x"05841188",
  7542 => x"150c8c08",
  7543 => x"ffa40508",
  7544 => x"8c08fcf4",
  7545 => x"050c5158",
  7546 => x"5858800b",
  7547 => x"8c08fcf0",
  7548 => x"050c8c08",
  7549 => x"ffac0508",
  7550 => x"8c08ffa8",
  7551 => x"05085757",
  7552 => x"84170884",
  7553 => x"17082e89",
  7554 => x"38810b8c",
  7555 => x"08fcf005",
  7556 => x"0c8c08fc",
  7557 => x"f405088c",
  7558 => x"08fcf005",
  7559 => x"0884120c",
  7560 => x"578c08ff",
  7561 => x"900508f8",
  7562 => x"0a268438",
  7563 => x"81a8398c",
  7564 => x"08ffa405",
  7565 => x"08881108",
  7566 => x"81058812",
  7567 => x"0c8c08ff",
  7568 => x"90050880",
  7569 => x"068c08ff",
  7570 => x"94050881",
  7571 => x"06705259",
  7572 => x"51567580",
  7573 => x"2e80cf38",
  7574 => x"8c08ff98",
  7575 => x"05089f2b",
  7576 => x"8c08ff9c",
  7577 => x"0508812a",
  7578 => x"7072078c",
  7579 => x"08ff9805",
  7580 => x"08812a59",
  7581 => x"59595975",
  7582 => x"8c08ff98",
  7583 => x"050c768c",
  7584 => x"08ff9c05",
  7585 => x"0c8c08ff",
  7586 => x"98050881",
  7587 => x"0a078c08",
  7588 => x"ff9c0508",
  7589 => x"80075856",
  7590 => x"758c08ff",
  7591 => x"98050c76",
  7592 => x"8c08ff9c",
  7593 => x"050c8c08",
  7594 => x"ff900508",
  7595 => x"9f2b8c08",
  7596 => x"ff940508",
  7597 => x"812a7072",
  7598 => x"078c08ff",
  7599 => x"90050881",
  7600 => x"2a595959",
  7601 => x"59758c08",
  7602 => x"ff90050c",
  7603 => x"768c08ff",
  7604 => x"94050cfe",
  7605 => x"cc398c08",
  7606 => x"ff900508",
  7607 => x"f00a2681",
  7608 => x"96388c08",
  7609 => x"ffa40508",
  7610 => x"881108ff",
  7611 => x"0588120c",
  7612 => x"8c08ff94",
  7613 => x"05089f2a",
  7614 => x"8c08ff90",
  7615 => x"05081070",
  7616 => x"72078c08",
  7617 => x"ff940508",
  7618 => x"105b535a",
  7619 => x"5a56758c",
  7620 => x"08ff9005",
  7621 => x"0c768c08",
  7622 => x"ff94050c",
  7623 => x"800b8c08",
  7624 => x"ff980508",
  7625 => x"248338a1",
  7626 => x"398c08ff",
  7627 => x"90050880",
  7628 => x"078c08ff",
  7629 => x"94050881",
  7630 => x"07585675",
  7631 => x"8c08ff90",
  7632 => x"050c768c",
  7633 => x"08ff9405",
  7634 => x"0c8c08ff",
  7635 => x"9c05089f",
  7636 => x"2a8c08ff",
  7637 => x"98050810",
  7638 => x"7072078c",
  7639 => x"08ff9c05",
  7640 => x"08105a58",
  7641 => x"5959758c",
  7642 => x"08ff9805",
  7643 => x"0c768c08",
  7644 => x"ff9c050c",
  7645 => x"fee0398c",
  7646 => x"08ff9005",
  7647 => x"08800670",
  7648 => x"8c08fce8",
  7649 => x"050c8c08",
  7650 => x"ff940508",
  7651 => x"81ff0670",
  7652 => x"8c08fcec",
  7653 => x"050c5856",
  7654 => x"8c08fce8",
  7655 => x"05088c08",
  7656 => x"fcec0508",
  7657 => x"5856758c",
  7658 => x"08fce805",
  7659 => x"0c768c08",
  7660 => x"fcec050c",
  7661 => x"8c08fce8",
  7662 => x"05085776",
  7663 => x"83bc388c",
  7664 => x"08fcec05",
  7665 => x"08567581",
  7666 => x"802e0981",
  7667 => x"0683ab38",
  7668 => x"8c08ff90",
  7669 => x"0508982b",
  7670 => x"8c08ff94",
  7671 => x"0508882a",
  7672 => x"7072078c",
  7673 => x"08ff9005",
  7674 => x"08882a71",
  7675 => x"81065159",
  7676 => x"59595975",
  7677 => x"802e81b8",
  7678 => x"388c08ff",
  7679 => x"9005088c",
  7680 => x"08ff9405",
  7681 => x"08585675",
  7682 => x"8c08fce0",
  7683 => x"050c768c",
  7684 => x"08fce405",
  7685 => x"0c805681",
  7686 => x"8057758c",
  7687 => x"08fcd805",
  7688 => x"0c768c08",
  7689 => x"fcdc050c",
  7690 => x"8c08fce4",
  7691 => x"05088c08",
  7692 => x"fcdc0508",
  7693 => x"7012708c",
  7694 => x"08fcd405",
  7695 => x"0c525757",
  7696 => x"810b8c08",
  7697 => x"fccc050c",
  7698 => x"8c08fcd4",
  7699 => x"05088c08",
  7700 => x"fce40508",
  7701 => x"57577577",
  7702 => x"26893880",
  7703 => x"0b8c08fc",
  7704 => x"cc050c8c",
  7705 => x"08fce005",
  7706 => x"088c08fc",
  7707 => x"d8050870",
  7708 => x"12708c08",
  7709 => x"fcd0050c",
  7710 => x"8c08fcd0",
  7711 => x"05088c08",
  7712 => x"fccc0508",
  7713 => x"11708c08",
  7714 => x"fcd0050c",
  7715 => x"53515257",
  7716 => x"578c08fc",
  7717 => x"d005088c",
  7718 => x"08fcd405",
  7719 => x"08585675",
  7720 => x"8c08ff90",
  7721 => x"050c768c",
  7722 => x"08ff9405",
  7723 => x"0c81cb39",
  7724 => x"8c08ff98",
  7725 => x"0508708c",
  7726 => x"08ff9c05",
  7727 => x"08075156",
  7728 => x"75802e81",
  7729 => x"b5388c08",
  7730 => x"ff900508",
  7731 => x"8c08ff94",
  7732 => x"05085856",
  7733 => x"758c08fc",
  7734 => x"c4050c76",
  7735 => x"8c08fcc8",
  7736 => x"050c8056",
  7737 => x"81805775",
  7738 => x"8c08fcbc",
  7739 => x"050c768c",
  7740 => x"08fcc005",
  7741 => x"0c8c08fc",
  7742 => x"c805088c",
  7743 => x"08fcc005",
  7744 => x"08701270",
  7745 => x"8c08fcb8",
  7746 => x"050c5257",
  7747 => x"57810b8c",
  7748 => x"08fcb005",
  7749 => x"0c8c08fc",
  7750 => x"b805088c",
  7751 => x"08fcc805",
  7752 => x"08575775",
  7753 => x"77268938",
  7754 => x"800b8c08",
  7755 => x"fcb0050c",
  7756 => x"8c08fcc4",
  7757 => x"05088c08",
  7758 => x"fcbc0508",
  7759 => x"7012708c",
  7760 => x"08fcb405",
  7761 => x"0c8c08fc",
  7762 => x"b405088c",
  7763 => x"08fcb005",
  7764 => x"0811708c",
  7765 => x"08fcb405",
  7766 => x"0c535152",
  7767 => x"57578c08",
  7768 => x"fcb40508",
  7769 => x"8c08fcb8",
  7770 => x"05085856",
  7771 => x"758c08ff",
  7772 => x"90050c76",
  7773 => x"8c08ff94",
  7774 => x"050c8c08",
  7775 => x"ffa40508",
  7776 => x"568c08ff",
  7777 => x"9005088c",
  7778 => x"08ff9405",
  7779 => x"08595776",
  7780 => x"8c170c77",
  7781 => x"90170c8c",
  7782 => x"08ffa405",
  7783 => x"08568376",
  7784 => x"0c8c08ff",
  7785 => x"a405088c",
  7786 => x"08ffa005",
  7787 => x"0c8c08ff",
  7788 => x"a0050870",
  7789 => x"8c08c005",
  7790 => x"0c8c08c0",
  7791 => x"0508538c",
  7792 => x"08880508",
  7793 => x"5256a8d0",
  7794 => x"3f8c0888",
  7795 => x"0508800c",
  7796 => x"80ff3d0d",
  7797 => x"8c0c048c",
  7798 => x"08028c0c",
  7799 => x"803d0d82",
  7800 => x"c08c7080",
  7801 => x"0c51823d",
  7802 => x"0d8c0c04",
  7803 => x"8c08028c",
  7804 => x"0cff3d0d",
  7805 => x"800b8c08",
  7806 => x"fc050c8c",
  7807 => x"08880508",
  7808 => x"51700882",
  7809 => x"2e098106",
  7810 => x"8838810b",
  7811 => x"8c08fc05",
  7812 => x"0c8c08fc",
  7813 => x"05087080",
  7814 => x"0c51833d",
  7815 => x"0d8c0c04",
  7816 => x"8c08028c",
  7817 => x"0cff3d0d",
  7818 => x"800b8c08",
  7819 => x"fc050c8c",
  7820 => x"08880508",
  7821 => x"51700884",
  7822 => x"2e098106",
  7823 => x"8838810b",
  7824 => x"8c08fc05",
  7825 => x"0c8c08fc",
  7826 => x"05087080",
  7827 => x"0c51833d",
  7828 => x"0d8c0c04",
  7829 => x"8c08028c",
  7830 => x"0cff3d0d",
  7831 => x"800b8c08",
  7832 => x"fc050c8c",
  7833 => x"08880508",
  7834 => x"51700880",
  7835 => x"2e8f388c",
  7836 => x"08880508",
  7837 => x"51700881",
  7838 => x"2e833888",
  7839 => x"39810b8c",
  7840 => x"08fc050c",
  7841 => x"8c08fc05",
  7842 => x"0870800c",
  7843 => x"51833d0d",
  7844 => x"8c0c048c",
  7845 => x"08028c0c",
  7846 => x"ffbc3d0d",
  7847 => x"8c088c05",
  7848 => x"088c0890",
  7849 => x"05085553",
  7850 => x"728c08cc",
  7851 => x"050c738c",
  7852 => x"08d0050c",
  7853 => x"8c089405",
  7854 => x"088c0898",
  7855 => x"05085553",
  7856 => x"728c08c4",
  7857 => x"050c738c",
  7858 => x"08c8050c",
  7859 => x"8c08ec05",
  7860 => x"70538c08",
  7861 => x"cc057053",
  7862 => x"5153b6f2",
  7863 => x"3f8c08d8",
  7864 => x"0570538c",
  7865 => x"08c40570",
  7866 => x"535153b6",
  7867 => x"e13f8c08",
  7868 => x"ec058c08",
  7869 => x"c0050c8c",
  7870 => x"08d8058c",
  7871 => x"08ffbc05",
  7872 => x"0c8c08c0",
  7873 => x"0508518e",
  7874 => x"fa3f8008",
  7875 => x"5372802e",
  7876 => x"8f388c08",
  7877 => x"c005088c",
  7878 => x"08ffb805",
  7879 => x"0c8dbd39",
  7880 => x"8c08ffbc",
  7881 => x"0508518e",
  7882 => x"da3f8008",
  7883 => x"5372802e",
  7884 => x"90388c08",
  7885 => x"ffbc0508",
  7886 => x"8c08ffb8",
  7887 => x"050c8d9c",
  7888 => x"398c08c0",
  7889 => x"05088c08",
  7890 => x"c005088c",
  7891 => x"08ffbc05",
  7892 => x"08841208",
  7893 => x"84120832",
  7894 => x"84140c8c",
  7895 => x"08c00508",
  7896 => x"54555555",
  7897 => x"8de93f80",
  7898 => x"08537292",
  7899 => x"388c08c0",
  7900 => x"0508518d",
  7901 => x"a63f8008",
  7902 => x"53728338",
  7903 => x"b6398c08",
  7904 => x"c005088c",
  7905 => x"08ffbc05",
  7906 => x"08545473",
  7907 => x"0873082e",
  7908 => x"09810691",
  7909 => x"388cef3f",
  7910 => x"8008708c",
  7911 => x"08ffb805",
  7912 => x"0c538cb8",
  7913 => x"398c08c0",
  7914 => x"05088c08",
  7915 => x"ffb8050c",
  7916 => x"8caa398c",
  7917 => x"08ffbc05",
  7918 => x"08518d93",
  7919 => x"3f800853",
  7920 => x"72802eac",
  7921 => x"388c08c0",
  7922 => x"05085380",
  7923 => x"54805573",
  7924 => x"8c140c74",
  7925 => x"90140c8c",
  7926 => x"08c00508",
  7927 => x"53800b88",
  7928 => x"140c8c08",
  7929 => x"c005088c",
  7930 => x"08ffb805",
  7931 => x"0c8bed39",
  7932 => x"8c08ffbc",
  7933 => x"0508518c",
  7934 => x"a23f8008",
  7935 => x"5372802e",
  7936 => x"98388c08",
  7937 => x"c0050853",
  7938 => x"84730c8c",
  7939 => x"08c00508",
  7940 => x"8c08ffb8",
  7941 => x"050c8bc4",
  7942 => x"398c08c0",
  7943 => x"05088c08",
  7944 => x"c005088c",
  7945 => x"08ffbc05",
  7946 => x"08881208",
  7947 => x"88120831",
  7948 => x"88140c8c",
  7949 => x"08c00508",
  7950 => x"51555555",
  7951 => x"9013088c",
  7952 => x"14085454",
  7953 => x"728c08ff",
  7954 => x"a8050c73",
  7955 => x"8c08ffac",
  7956 => x"050c8c08",
  7957 => x"ffbc0508",
  7958 => x"53901308",
  7959 => x"8c140854",
  7960 => x"54728c08",
  7961 => x"ffa0050c",
  7962 => x"738c08ff",
  7963 => x"a4050c8c",
  7964 => x"08ffa005",
  7965 => x"088c08ff",
  7966 => x"a8050826",
  7967 => x"a6388c08",
  7968 => x"ffa00508",
  7969 => x"8c08ffa8",
  7970 => x"05082e09",
  7971 => x"810681de",
  7972 => x"388c08ff",
  7973 => x"a405088c",
  7974 => x"08ffac05",
  7975 => x"08268438",
  7976 => x"81cc398c",
  7977 => x"08ffa805",
  7978 => x"088c08ff",
  7979 => x"ac050855",
  7980 => x"53728c08",
  7981 => x"ff90050c",
  7982 => x"738c08ff",
  7983 => x"94050c8c",
  7984 => x"08ff9005",
  7985 => x"088c08ff",
  7986 => x"94050855",
  7987 => x"53728c08",
  7988 => x"ff88050c",
  7989 => x"738c08ff",
  7990 => x"8c050c8c",
  7991 => x"08ff8c05",
  7992 => x"088c08ff",
  7993 => x"94050870",
  7994 => x"12708c08",
  7995 => x"ff84050c",
  7996 => x"52545481",
  7997 => x"0b8c08fe",
  7998 => x"fc050c8c",
  7999 => x"08ff8405",
  8000 => x"088c08ff",
  8001 => x"8c050854",
  8002 => x"54727426",
  8003 => x"8938800b",
  8004 => x"8c08fefc",
  8005 => x"050c8c08",
  8006 => x"ff880508",
  8007 => x"8c08ff90",
  8008 => x"05087012",
  8009 => x"708c08ff",
  8010 => x"80050c8c",
  8011 => x"08ff8005",
  8012 => x"088c08fe",
  8013 => x"fc050811",
  8014 => x"708c08ff",
  8015 => x"80050c53",
  8016 => x"51525454",
  8017 => x"8c08ff80",
  8018 => x"05088c08",
  8019 => x"ff840508",
  8020 => x"5553728c",
  8021 => x"08ffa805",
  8022 => x"0c738c08",
  8023 => x"ffac050c",
  8024 => x"8c08c005",
  8025 => x"08881108",
  8026 => x"ff058812",
  8027 => x"0c53880a",
  8028 => x"53805472",
  8029 => x"8c08ffb0",
  8030 => x"050c738c",
  8031 => x"08ffb405",
  8032 => x"0c805380",
  8033 => x"54728c08",
  8034 => x"ff98050c",
  8035 => x"738c08ff",
  8036 => x"9c050c8c",
  8037 => x"08ffb005",
  8038 => x"08708c08",
  8039 => x"ffb40508",
  8040 => x"07515372",
  8041 => x"802e848a",
  8042 => x"388c08ff",
  8043 => x"a005088c",
  8044 => x"08ffa805",
  8045 => x"0826828d",
  8046 => x"388c08ff",
  8047 => x"a005088c",
  8048 => x"08ffa805",
  8049 => x"082e0981",
  8050 => x"0691388c",
  8051 => x"08ffa405",
  8052 => x"088c08ff",
  8053 => x"ac050826",
  8054 => x"81eb388c",
  8055 => x"08ff9805",
  8056 => x"088c08ff",
  8057 => x"b0050807",
  8058 => x"8c08ff9c",
  8059 => x"05088c08",
  8060 => x"ffb40508",
  8061 => x"07555372",
  8062 => x"8c08ff98",
  8063 => x"050c738c",
  8064 => x"08ff9c05",
  8065 => x"0c8c08ff",
  8066 => x"a805088c",
  8067 => x"08ffac05",
  8068 => x"08555372",
  8069 => x"8c08fef4",
  8070 => x"050c738c",
  8071 => x"08fef805",
  8072 => x"0c8c08ff",
  8073 => x"a005088c",
  8074 => x"08ffa405",
  8075 => x"08555372",
  8076 => x"8c08feec",
  8077 => x"050c738c",
  8078 => x"08fef005",
  8079 => x"0c8c08fe",
  8080 => x"f805088c",
  8081 => x"08fef005",
  8082 => x"08717131",
  8083 => x"708c08fe",
  8084 => x"e8050c52",
  8085 => x"5454810b",
  8086 => x"8c08fee0",
  8087 => x"050c8c08",
  8088 => x"fee80508",
  8089 => x"8c08fef8",
  8090 => x"05085454",
  8091 => x"73732689",
  8092 => x"38800b8c",
  8093 => x"08fee005",
  8094 => x"0c8c08fe",
  8095 => x"f405088c",
  8096 => x"08feec05",
  8097 => x"08717131",
  8098 => x"708c08fe",
  8099 => x"e4050c8c",
  8100 => x"08fee405",
  8101 => x"08708c08",
  8102 => x"fee00508",
  8103 => x"31708c08",
  8104 => x"fee4050c",
  8105 => x"53515254",
  8106 => x"548c08fe",
  8107 => x"e405088c",
  8108 => x"08fee805",
  8109 => x"08555372",
  8110 => x"8c08ffa8",
  8111 => x"050c738c",
  8112 => x"08ffac05",
  8113 => x"0c8c08ff",
  8114 => x"b005089f",
  8115 => x"2b8c08ff",
  8116 => x"b4050881",
  8117 => x"2a707207",
  8118 => x"8c08ffb0",
  8119 => x"0508812a",
  8120 => x"56565656",
  8121 => x"728c08ff",
  8122 => x"b0050c73",
  8123 => x"8c08ffb4",
  8124 => x"050c8c08",
  8125 => x"ffa80508",
  8126 => x"8c08ffac",
  8127 => x"05085553",
  8128 => x"728c08fe",
  8129 => x"d8050c73",
  8130 => x"8c08fedc",
  8131 => x"050c8c08",
  8132 => x"fed80508",
  8133 => x"8c08fedc",
  8134 => x"05085553",
  8135 => x"728c08fe",
  8136 => x"d0050c73",
  8137 => x"8c08fed4",
  8138 => x"050c8c08",
  8139 => x"fed40508",
  8140 => x"8c08fedc",
  8141 => x"05087012",
  8142 => x"708c08fe",
  8143 => x"cc050c52",
  8144 => x"5454810b",
  8145 => x"8c08fec4",
  8146 => x"050c8c08",
  8147 => x"fecc0508",
  8148 => x"8c08fed4",
  8149 => x"05085454",
  8150 => x"72742689",
  8151 => x"38800b8c",
  8152 => x"08fec405",
  8153 => x"0c8c08fe",
  8154 => x"d005088c",
  8155 => x"08fed805",
  8156 => x"08701270",
  8157 => x"8c08fec8",
  8158 => x"050c8c08",
  8159 => x"fec80508",
  8160 => x"8c08fec4",
  8161 => x"05081170",
  8162 => x"8c08fec8",
  8163 => x"050c5351",
  8164 => x"5254548c",
  8165 => x"08fec805",
  8166 => x"088c08fe",
  8167 => x"cc050855",
  8168 => x"53728c08",
  8169 => x"ffa8050c",
  8170 => x"738c08ff",
  8171 => x"ac050cfb",
  8172 => x"e2398c08",
  8173 => x"ff980508",
  8174 => x"8006708c",
  8175 => x"08febc05",
  8176 => x"0c8c08ff",
  8177 => x"9c050881",
  8178 => x"ff06708c",
  8179 => x"08fec005",
  8180 => x"0c54548c",
  8181 => x"08febc05",
  8182 => x"088c08fe",
  8183 => x"c0050855",
  8184 => x"53728c08",
  8185 => x"febc050c",
  8186 => x"738c08fe",
  8187 => x"c0050c8c",
  8188 => x"08febc05",
  8189 => x"08547383",
  8190 => x"bc388c08",
  8191 => x"fec00508",
  8192 => x"53728180",
  8193 => x"2e098106",
  8194 => x"83ab388c",
  8195 => x"08ff9805",
  8196 => x"08982b8c",
  8197 => x"08ff9c05",
  8198 => x"08882a70",
  8199 => x"72078c08",
  8200 => x"ff980508",
  8201 => x"882a7181",
  8202 => x"06515656",
  8203 => x"56567280",
  8204 => x"2e81b838",
  8205 => x"8c08ff98",
  8206 => x"05088c08",
  8207 => x"ff9c0508",
  8208 => x"5553728c",
  8209 => x"08feb405",
  8210 => x"0c738c08",
  8211 => x"feb8050c",
  8212 => x"80538180",
  8213 => x"54728c08",
  8214 => x"feac050c",
  8215 => x"738c08fe",
  8216 => x"b0050c8c",
  8217 => x"08feb805",
  8218 => x"088c08fe",
  8219 => x"b0050870",
  8220 => x"12708c08",
  8221 => x"fea8050c",
  8222 => x"52545481",
  8223 => x"0b8c08fe",
  8224 => x"a0050c8c",
  8225 => x"08fea805",
  8226 => x"088c08fe",
  8227 => x"b8050854",
  8228 => x"54727426",
  8229 => x"8938800b",
  8230 => x"8c08fea0",
  8231 => x"050c8c08",
  8232 => x"feb40508",
  8233 => x"8c08feac",
  8234 => x"05087012",
  8235 => x"708c08fe",
  8236 => x"a4050c8c",
  8237 => x"08fea405",
  8238 => x"088c08fe",
  8239 => x"a0050811",
  8240 => x"708c08fe",
  8241 => x"a4050c53",
  8242 => x"51525454",
  8243 => x"8c08fea4",
  8244 => x"05088c08",
  8245 => x"fea80508",
  8246 => x"5553728c",
  8247 => x"08ff9805",
  8248 => x"0c738c08",
  8249 => x"ff9c050c",
  8250 => x"81cb398c",
  8251 => x"08ffa805",
  8252 => x"08708c08",
  8253 => x"ffac0508",
  8254 => x"07515372",
  8255 => x"802e81b5",
  8256 => x"388c08ff",
  8257 => x"9805088c",
  8258 => x"08ff9c05",
  8259 => x"08555372",
  8260 => x"8c08fe98",
  8261 => x"050c738c",
  8262 => x"08fe9c05",
  8263 => x"0c805381",
  8264 => x"8054728c",
  8265 => x"08fe9005",
  8266 => x"0c738c08",
  8267 => x"fe94050c",
  8268 => x"8c08fe9c",
  8269 => x"05088c08",
  8270 => x"fe940508",
  8271 => x"7012708c",
  8272 => x"08fe8c05",
  8273 => x"0c525454",
  8274 => x"810b8c08",
  8275 => x"fe84050c",
  8276 => x"8c08fe8c",
  8277 => x"05088c08",
  8278 => x"fe9c0508",
  8279 => x"54547274",
  8280 => x"26893880",
  8281 => x"0b8c08fe",
  8282 => x"84050c8c",
  8283 => x"08fe9805",
  8284 => x"088c08fe",
  8285 => x"90050870",
  8286 => x"12708c08",
  8287 => x"fe88050c",
  8288 => x"8c08fe88",
  8289 => x"05088c08",
  8290 => x"fe840508",
  8291 => x"11708c08",
  8292 => x"fe88050c",
  8293 => x"53515254",
  8294 => x"548c08fe",
  8295 => x"8805088c",
  8296 => x"08fe8c05",
  8297 => x"08555372",
  8298 => x"8c08ff98",
  8299 => x"050c738c",
  8300 => x"08ff9c05",
  8301 => x"0c8c08c0",
  8302 => x"0508558c",
  8303 => x"08ff9805",
  8304 => x"088c08ff",
  8305 => x"9c050855",
  8306 => x"53728c16",
  8307 => x"0c739016",
  8308 => x"0c8c08c0",
  8309 => x"05088c08",
  8310 => x"ffb8050c",
  8311 => x"8c08ffb8",
  8312 => x"0508708c",
  8313 => x"08d4050c",
  8314 => x"8c08d405",
  8315 => x"08538c08",
  8316 => x"88050852",
  8317 => x"5398a13f",
  8318 => x"8c088805",
  8319 => x"08800c80",
  8320 => x"c63d0d8c",
  8321 => x"0c048c08",
  8322 => x"028c0c80",
  8323 => x"3d0d82c0",
  8324 => x"8c70800c",
  8325 => x"51823d0d",
  8326 => x"8c0c048c",
  8327 => x"08028c0c",
  8328 => x"ff3d0d80",
  8329 => x"0b8c08fc",
  8330 => x"050c8c08",
  8331 => x"88050851",
  8332 => x"7008822e",
  8333 => x"09810688",
  8334 => x"38810b8c",
  8335 => x"08fc050c",
  8336 => x"8c08fc05",
  8337 => x"0870800c",
  8338 => x"51833d0d",
  8339 => x"8c0c048c",
  8340 => x"08028c0c",
  8341 => x"ff3d0d80",
  8342 => x"0b8c08fc",
  8343 => x"050c8c08",
  8344 => x"88050851",
  8345 => x"7008842e",
  8346 => x"09810688",
  8347 => x"38810b8c",
  8348 => x"08fc050c",
  8349 => x"8c08fc05",
  8350 => x"0870800c",
  8351 => x"51833d0d",
  8352 => x"8c0c048c",
  8353 => x"08028c0c",
  8354 => x"ff3d0d80",
  8355 => x"0b8c08fc",
  8356 => x"050c8c08",
  8357 => x"88050851",
  8358 => x"7008802e",
  8359 => x"8f388c08",
  8360 => x"88050851",
  8361 => x"7008812e",
  8362 => x"83388839",
  8363 => x"810b8c08",
  8364 => x"fc050c8c",
  8365 => x"08fc0508",
  8366 => x"70800c51",
  8367 => x"833d0d8c",
  8368 => x"0c048c08",
  8369 => x"028c0cee",
  8370 => x"3d0d8c08",
  8371 => x"8805088c",
  8372 => x"088c0508",
  8373 => x"5553728c",
  8374 => x"08d0050c",
  8375 => x"738c08d4",
  8376 => x"050c8c08",
  8377 => x"9005088c",
  8378 => x"08940508",
  8379 => x"5553728c",
  8380 => x"08c8050c",
  8381 => x"738c08cc",
  8382 => x"050c8c08",
  8383 => x"ec057053",
  8384 => x"8c08d005",
  8385 => x"70535153",
  8386 => x"a6c43f8c",
  8387 => x"08d80570",
  8388 => x"538c08c8",
  8389 => x"05705351",
  8390 => x"53a6b33f",
  8391 => x"8c08ec05",
  8392 => x"70525380",
  8393 => x"c83f8008",
  8394 => x"53729238",
  8395 => x"8c08d805",
  8396 => x"705253b9",
  8397 => x"3f800853",
  8398 => x"7283388a",
  8399 => x"39810b8c",
  8400 => x"08c4050c",
  8401 => x"9b398c08",
  8402 => x"d8057053",
  8403 => x"8c08ec05",
  8404 => x"70535153",
  8405 => x"a9d63f80",
  8406 => x"08708c08",
  8407 => x"c4050c53",
  8408 => x"8c08c405",
  8409 => x"08800c94",
  8410 => x"3d0d8c0c",
  8411 => x"048c0802",
  8412 => x"8c0cff3d",
  8413 => x"0d800b8c",
  8414 => x"08fc050c",
  8415 => x"8c088805",
  8416 => x"08517008",
  8417 => x"802e8f38",
  8418 => x"8c088805",
  8419 => x"08517008",
  8420 => x"812e8338",
  8421 => x"8839810b",
  8422 => x"8c08fc05",
  8423 => x"0c8c08fc",
  8424 => x"05087080",
  8425 => x"0c51833d",
  8426 => x"0d8c0c04",
  8427 => x"8c08028c",
  8428 => x"0cee3d0d",
  8429 => x"8c088805",
  8430 => x"088c088c",
  8431 => x"05085553",
  8432 => x"728c08d0",
  8433 => x"050c738c",
  8434 => x"08d4050c",
  8435 => x"8c089005",
  8436 => x"088c0894",
  8437 => x"05085553",
  8438 => x"728c08c8",
  8439 => x"050c738c",
  8440 => x"08cc050c",
  8441 => x"8c08ec05",
  8442 => x"70538c08",
  8443 => x"d0057053",
  8444 => x"5153a4da",
  8445 => x"3f8c08d8",
  8446 => x"0570538c",
  8447 => x"08c80570",
  8448 => x"535153a4",
  8449 => x"c93f8c08",
  8450 => x"ec057052",
  8451 => x"5380c83f",
  8452 => x"80085372",
  8453 => x"92388c08",
  8454 => x"d8057052",
  8455 => x"53b93f80",
  8456 => x"08537283",
  8457 => x"388a3981",
  8458 => x"0b8c08c4",
  8459 => x"050c9b39",
  8460 => x"8c08d805",
  8461 => x"70538c08",
  8462 => x"ec057053",
  8463 => x"5153a7ec",
  8464 => x"3f800870",
  8465 => x"8c08c405",
  8466 => x"0c538c08",
  8467 => x"c4050880",
  8468 => x"0c943d0d",
  8469 => x"8c0c048c",
  8470 => x"08028c0c",
  8471 => x"ff3d0d80",
  8472 => x"0b8c08fc",
  8473 => x"050c8c08",
  8474 => x"88050851",
  8475 => x"7008802e",
  8476 => x"8f388c08",
  8477 => x"88050851",
  8478 => x"7008812e",
  8479 => x"83388839",
  8480 => x"810b8c08",
  8481 => x"fc050c8c",
  8482 => x"08fc0508",
  8483 => x"70800c51",
  8484 => x"833d0d8c",
  8485 => x"0c048c08",
  8486 => x"028c0cee",
  8487 => x"3d0d8c08",
  8488 => x"8805088c",
  8489 => x"088c0508",
  8490 => x"5553728c",
  8491 => x"08d0050c",
  8492 => x"738c08d4",
  8493 => x"050c8c08",
  8494 => x"9005088c",
  8495 => x"08940508",
  8496 => x"5553728c",
  8497 => x"08c8050c",
  8498 => x"738c08cc",
  8499 => x"050c8c08",
  8500 => x"ec057053",
  8501 => x"8c08d005",
  8502 => x"70535153",
  8503 => x"a2f03f8c",
  8504 => x"08d80570",
  8505 => x"538c08c8",
  8506 => x"05705351",
  8507 => x"53a2df3f",
  8508 => x"8c08ec05",
  8509 => x"70525380",
  8510 => x"c83f8008",
  8511 => x"53729238",
  8512 => x"8c08d805",
  8513 => x"705253b9",
  8514 => x"3f800853",
  8515 => x"7283388a",
  8516 => x"39ff0b8c",
  8517 => x"08c4050c",
  8518 => x"9b398c08",
  8519 => x"d8057053",
  8520 => x"8c08ec05",
  8521 => x"70535153",
  8522 => x"a6823f80",
  8523 => x"08708c08",
  8524 => x"c4050c53",
  8525 => x"8c08c405",
  8526 => x"08800c94",
  8527 => x"3d0d8c0c",
  8528 => x"048c0802",
  8529 => x"8c0cff3d",
  8530 => x"0d800b8c",
  8531 => x"08fc050c",
  8532 => x"8c088805",
  8533 => x"08517008",
  8534 => x"802e8f38",
  8535 => x"8c088805",
  8536 => x"08517008",
  8537 => x"812e8338",
  8538 => x"8839810b",
  8539 => x"8c08fc05",
  8540 => x"0c8c08fc",
  8541 => x"05087080",
  8542 => x"0c51833d",
  8543 => x"0d8c0c04",
  8544 => x"8c08028c",
  8545 => x"0cee3d0d",
  8546 => x"8c088805",
  8547 => x"088c088c",
  8548 => x"05085553",
  8549 => x"728c08d0",
  8550 => x"050c738c",
  8551 => x"08d4050c",
  8552 => x"8c089005",
  8553 => x"088c0894",
  8554 => x"05085553",
  8555 => x"728c08c8",
  8556 => x"050c738c",
  8557 => x"08cc050c",
  8558 => x"8c08ec05",
  8559 => x"70538c08",
  8560 => x"d0057053",
  8561 => x"5153a186",
  8562 => x"3f8c08d8",
  8563 => x"0570538c",
  8564 => x"08c80570",
  8565 => x"535153a0",
  8566 => x"f53f8c08",
  8567 => x"ec057052",
  8568 => x"5380c83f",
  8569 => x"80085372",
  8570 => x"92388c08",
  8571 => x"d8057052",
  8572 => x"53b93f80",
  8573 => x"08537283",
  8574 => x"388a3981",
  8575 => x"0b8c08c4",
  8576 => x"050c9b39",
  8577 => x"8c08d805",
  8578 => x"70538c08",
  8579 => x"ec057053",
  8580 => x"5153a498",
  8581 => x"3f800870",
  8582 => x"8c08c405",
  8583 => x"0c538c08",
  8584 => x"c4050880",
  8585 => x"0c943d0d",
  8586 => x"8c0c048c",
  8587 => x"08028c0c",
  8588 => x"ff3d0d80",
  8589 => x"0b8c08fc",
  8590 => x"050c8c08",
  8591 => x"88050851",
  8592 => x"7008802e",
  8593 => x"8f388c08",
  8594 => x"88050851",
  8595 => x"7008812e",
  8596 => x"83388839",
  8597 => x"810b8c08",
  8598 => x"fc050c8c",
  8599 => x"08fc0508",
  8600 => x"70800c51",
  8601 => x"833d0d8c",
  8602 => x"0c048c08",
  8603 => x"028c0cee",
  8604 => x"3d0d8c08",
  8605 => x"8805088c",
  8606 => x"088c0508",
  8607 => x"5553728c",
  8608 => x"08d0050c",
  8609 => x"738c08d4",
  8610 => x"050c8c08",
  8611 => x"9005088c",
  8612 => x"08940508",
  8613 => x"5553728c",
  8614 => x"08c8050c",
  8615 => x"738c08cc",
  8616 => x"050c8c08",
  8617 => x"ec057053",
  8618 => x"8c08d005",
  8619 => x"70535153",
  8620 => x"9f9c3f8c",
  8621 => x"08d80570",
  8622 => x"538c08c8",
  8623 => x"05705351",
  8624 => x"539f8b3f",
  8625 => x"8c08ec05",
  8626 => x"70525380",
  8627 => x"c83f8008",
  8628 => x"53729238",
  8629 => x"8c08d805",
  8630 => x"705253b9",
  8631 => x"3f800853",
  8632 => x"7283388a",
  8633 => x"39810b8c",
  8634 => x"08c4050c",
  8635 => x"9b398c08",
  8636 => x"d8057053",
  8637 => x"8c08ec05",
  8638 => x"70535153",
  8639 => x"a2ae3f80",
  8640 => x"08708c08",
  8641 => x"c4050c53",
  8642 => x"8c08c405",
  8643 => x"08800c94",
  8644 => x"3d0d8c0c",
  8645 => x"048c0802",
  8646 => x"8c0cff3d",
  8647 => x"0d800b8c",
  8648 => x"08fc050c",
  8649 => x"8c088805",
  8650 => x"08517008",
  8651 => x"802e8f38",
  8652 => x"8c088805",
  8653 => x"08517008",
  8654 => x"812e8338",
  8655 => x"8839810b",
  8656 => x"8c08fc05",
  8657 => x"0c8c08fc",
  8658 => x"05087080",
  8659 => x"0c51833d",
  8660 => x"0d8c0c04",
  8661 => x"8c08028c",
  8662 => x"0cf63d0d",
  8663 => x"830b8c08",
  8664 => x"ec050c80",
  8665 => x"0b8c08e8",
  8666 => x"050c8c08",
  8667 => x"8c050880",
  8668 => x"25883881",
  8669 => x"0b8c08e8",
  8670 => x"050c8c08",
  8671 => x"e805088c",
  8672 => x"08f0050c",
  8673 => x"8c088c05",
  8674 => x"088b3882",
  8675 => x"0b8c08ec",
  8676 => x"050c819e",
  8677 => x"39bc0b8c",
  8678 => x"08f4050c",
  8679 => x"8c08f005",
  8680 => x"08802ebe",
  8681 => x"388c088c",
  8682 => x"0508810a",
  8683 => x"2e098106",
  8684 => x"98388f83",
  8685 => x"0a53800b",
  8686 => x"8c088805",
  8687 => x"08565472",
  8688 => x"750c7384",
  8689 => x"160c80fa",
  8690 => x"398c088c",
  8691 => x"05083070",
  8692 => x"8c08fc05",
  8693 => x"0c709f2c",
  8694 => x"708c08f8",
  8695 => x"050c5153",
  8696 => x"97398c08",
  8697 => x"8c050870",
  8698 => x"8c08fc05",
  8699 => x"0c709f2c",
  8700 => x"708c08f8",
  8701 => x"050c5153",
  8702 => x"8c08f805",
  8703 => x"08f00a26",
  8704 => x"b1388c08",
  8705 => x"fc05089f",
  8706 => x"2a8c08f8",
  8707 => x"05081070",
  8708 => x"72078c08",
  8709 => x"f8050c8c",
  8710 => x"08fc0508",
  8711 => x"108c08fc",
  8712 => x"050c8c08",
  8713 => x"f40508ff",
  8714 => x"058c08f4",
  8715 => x"050c5454",
  8716 => x"c7398c08",
  8717 => x"ec057053",
  8718 => x"8c088805",
  8719 => x"0852538b",
  8720 => x"d73f8c08",
  8721 => x"88050880",
  8722 => x"0c8c3d0d",
  8723 => x"8c0c048c",
  8724 => x"08028c0c",
  8725 => x"ec3d0d8c",
  8726 => x"08880508",
  8727 => x"8c088c05",
  8728 => x"08575574",
  8729 => x"8c08e005",
  8730 => x"0c758c08",
  8731 => x"e4050c8c",
  8732 => x"08ec0570",
  8733 => x"538c08e0",
  8734 => x"05705351",
  8735 => x"559bcf3f",
  8736 => x"8c08ec05",
  8737 => x"70525583",
  8738 => x"8d3f8008",
  8739 => x"5574802e",
  8740 => x"8b38800b",
  8741 => x"8c08d405",
  8742 => x"0c81fb39",
  8743 => x"8c08ec05",
  8744 => x"70525582",
  8745 => x"b23f8008",
  8746 => x"5574802e",
  8747 => x"8b38800b",
  8748 => x"8c08d405",
  8749 => x"0c81df39",
  8750 => x"8c08ec05",
  8751 => x"70525581",
  8752 => x"e23f8008",
  8753 => x"5574802e",
  8754 => x"a9388c08",
  8755 => x"f0050880",
  8756 => x"2e8b3881",
  8757 => x"0a0b8c08",
  8758 => x"d0050c89",
  8759 => x"39fe0a0b",
  8760 => x"8c08d005",
  8761 => x"0c8c08d0",
  8762 => x"05088c08",
  8763 => x"d4050c81",
  8764 => x"a5398c08",
  8765 => x"f4050880",
  8766 => x"258b3880",
  8767 => x"0b8c08d4",
  8768 => x"050c8192",
  8769 => x"399e0b8c",
  8770 => x"08f40508",
  8771 => x"25a9388c",
  8772 => x"08f00508",
  8773 => x"802e8b38",
  8774 => x"810a0b8c",
  8775 => x"08cc050c",
  8776 => x"8939fe0a",
  8777 => x"0b8c08cc",
  8778 => x"050c8c08",
  8779 => x"cc05088c",
  8780 => x"08d4050c",
  8781 => x"80e039bc",
  8782 => x"0b8c08f4",
  8783 => x"0508318c",
  8784 => x"08d80571",
  8785 => x"5658558c",
  8786 => x"08f80508",
  8787 => x"8c08fc05",
  8788 => x"08575574",
  8789 => x"52755376",
  8790 => x"5187c63f",
  8791 => x"8c08d805",
  8792 => x"088c08dc",
  8793 => x"0508708c",
  8794 => x"08e8050c",
  8795 => x"8c08e805",
  8796 => x"088c08c8",
  8797 => x"050c5755",
  8798 => x"8c08f005",
  8799 => x"08802e8c",
  8800 => x"388c08c8",
  8801 => x"0508308c",
  8802 => x"08c8050c",
  8803 => x"8c08c805",
  8804 => x"088c08d4",
  8805 => x"050c8c08",
  8806 => x"d4050880",
  8807 => x"0c963d0d",
  8808 => x"8c0c048c",
  8809 => x"08028c0c",
  8810 => x"ff3d0d80",
  8811 => x"0b8c08fc",
  8812 => x"050c8c08",
  8813 => x"88050851",
  8814 => x"7008842e",
  8815 => x"09810688",
  8816 => x"38810b8c",
  8817 => x"08fc050c",
  8818 => x"8c08fc05",
  8819 => x"0870800c",
  8820 => x"51833d0d",
  8821 => x"8c0c048c",
  8822 => x"08028c0c",
  8823 => x"ff3d0d80",
  8824 => x"0b8c08fc",
  8825 => x"050c8c08",
  8826 => x"88050851",
  8827 => x"7008802e",
  8828 => x"8f388c08",
  8829 => x"88050851",
  8830 => x"7008812e",
  8831 => x"83388839",
  8832 => x"810b8c08",
  8833 => x"fc050c8c",
  8834 => x"08fc0508",
  8835 => x"70800c51",
  8836 => x"833d0d8c",
  8837 => x"0c048c08",
  8838 => x"028c0cff",
  8839 => x"3d0d800b",
  8840 => x"8c08fc05",
  8841 => x"0c8c0888",
  8842 => x"05085170",
  8843 => x"08822e09",
  8844 => x"81068838",
  8845 => x"810b8c08",
  8846 => x"fc050c8c",
  8847 => x"08fc0508",
  8848 => x"70800c51",
  8849 => x"833d0d8c",
  8850 => x"0c048c08",
  8851 => x"028c0cfd",
  8852 => x"3d0d8053",
  8853 => x"8c088c05",
  8854 => x"08528c08",
  8855 => x"88050851",
  8856 => x"fdfba83f",
  8857 => x"80087080",
  8858 => x"0c54853d",
  8859 => x"0d8c0c04",
  8860 => x"8c08028c",
  8861 => x"0cfd3d0d",
  8862 => x"81538c08",
  8863 => x"8c050852",
  8864 => x"8c088805",
  8865 => x"0851fdfb",
  8866 => x"823f8008",
  8867 => x"70800c54",
  8868 => x"853d0d8c",
  8869 => x"0c048c08",
  8870 => x"028c0ceb",
  8871 => x"3d0d800b",
  8872 => x"8c08f005",
  8873 => x"0c800b8c",
  8874 => x"08f4050c",
  8875 => x"8c088c05",
  8876 => x"088c0890",
  8877 => x"05085654",
  8878 => x"738c08f0",
  8879 => x"050c748c",
  8880 => x"08f4050c",
  8881 => x"8c08f805",
  8882 => x"8c08f005",
  8883 => x"56568870",
  8884 => x"54755376",
  8885 => x"5254fdfc",
  8886 => x"b63f800b",
  8887 => x"8c08e805",
  8888 => x"0c800b8c",
  8889 => x"08ec050c",
  8890 => x"8c089405",
  8891 => x"088c0898",
  8892 => x"05085654",
  8893 => x"738c08e8",
  8894 => x"050c748c",
  8895 => x"08ec050c",
  8896 => x"8c08f005",
  8897 => x"8c08e805",
  8898 => x"56568870",
  8899 => x"54755376",
  8900 => x"5254fdfb",
  8901 => x"fa3f800b",
  8902 => x"8c08e805",
  8903 => x"0c800b8c",
  8904 => x"08ec050c",
  8905 => x"8c08fc05",
  8906 => x"0883ffff",
  8907 => x"068c08cc",
  8908 => x"050c8c08",
  8909 => x"fc050890",
  8910 => x"2a8c08c4",
  8911 => x"050c8c08",
  8912 => x"f4050883",
  8913 => x"ffff068c",
  8914 => x"08c8050c",
  8915 => x"8c08f405",
  8916 => x"08902a8c",
  8917 => x"08c0050c",
  8918 => x"8c08cc05",
  8919 => x"088c08c8",
  8920 => x"05082970",
  8921 => x"8c08dc05",
  8922 => x"0c8c08cc",
  8923 => x"05088c08",
  8924 => x"c0050829",
  8925 => x"708c08d8",
  8926 => x"050c8c08",
  8927 => x"c405088c",
  8928 => x"08c80508",
  8929 => x"29708c08",
  8930 => x"d4050c8c",
  8931 => x"08c40508",
  8932 => x"8c08c005",
  8933 => x"0829708c",
  8934 => x"08d0050c",
  8935 => x"8c08dc05",
  8936 => x"08902a8c",
  8937 => x"08d80508",
  8938 => x"118c08d8",
  8939 => x"050c8c08",
  8940 => x"d805088c",
  8941 => x"08d40508",
  8942 => x"058c08d8",
  8943 => x"050c5151",
  8944 => x"5151548c",
  8945 => x"08d80508",
  8946 => x"8c08d405",
  8947 => x"08278f38",
  8948 => x"8c08d005",
  8949 => x"08848080",
  8950 => x"058c08d0",
  8951 => x"050c8c08",
  8952 => x"d8050890",
  8953 => x"2a8c08d0",
  8954 => x"0508118c",
  8955 => x"08e0050c",
  8956 => x"8c08d805",
  8957 => x"0883ffff",
  8958 => x"0670902b",
  8959 => x"8c08dc05",
  8960 => x"0883ffff",
  8961 => x"0670128c",
  8962 => x"08e4050c",
  8963 => x"52575154",
  8964 => x"8c08e005",
  8965 => x"088c08e4",
  8966 => x"05085654",
  8967 => x"738c08e8",
  8968 => x"050c748c",
  8969 => x"08ec050c",
  8970 => x"8c08fc05",
  8971 => x"088c08f0",
  8972 => x"0508298c",
  8973 => x"08f80508",
  8974 => x"8c08f405",
  8975 => x"08297012",
  8976 => x"8c08e805",
  8977 => x"08118c08",
  8978 => x"e8050c51",
  8979 => x"55558c08",
  8980 => x"e805088c",
  8981 => x"08ec0508",
  8982 => x"8c088805",
  8983 => x"08585654",
  8984 => x"73760c74",
  8985 => x"84170c8c",
  8986 => x"08880508",
  8987 => x"800c973d",
  8988 => x"0d8c0c04",
  8989 => x"8c08028c",
  8990 => x"0cf63d0d",
  8991 => x"800b8c08",
  8992 => x"f0050c80",
  8993 => x"0b8c08f4",
  8994 => x"050c8c08",
  8995 => x"8c05088c",
  8996 => x"08900508",
  8997 => x"5654738c",
  8998 => x"08f0050c",
  8999 => x"748c08f4",
  9000 => x"050c8c08",
  9001 => x"f8058c08",
  9002 => x"f0055656",
  9003 => x"88705475",
  9004 => x"53765254",
  9005 => x"fdf8d83f",
  9006 => x"800b8c08",
  9007 => x"f0050c80",
  9008 => x"0b8c08f4",
  9009 => x"050c8c08",
  9010 => x"f8050830",
  9011 => x"8c08ec05",
  9012 => x"0c8c08fc",
  9013 => x"0508802e",
  9014 => x"8d388c08",
  9015 => x"ec0508ff",
  9016 => x"058c08ec",
  9017 => x"050c8c08",
  9018 => x"ec05088c",
  9019 => x"08f0050c",
  9020 => x"8c08fc05",
  9021 => x"08308c08",
  9022 => x"f4050c8c",
  9023 => x"08f00508",
  9024 => x"8c08f405",
  9025 => x"088c0888",
  9026 => x"05085856",
  9027 => x"5473760c",
  9028 => x"7484170c",
  9029 => x"8c088805",
  9030 => x"08800c8c",
  9031 => x"3d0d8c0c",
  9032 => x"048c0802",
  9033 => x"8c0cf53d",
  9034 => x"0d8c0894",
  9035 => x"05089d38",
  9036 => x"8c088c05",
  9037 => x"088c0890",
  9038 => x"05088c08",
  9039 => x"88050858",
  9040 => x"56547376",
  9041 => x"0c748417",
  9042 => x"0c81c039",
  9043 => x"800b8c08",
  9044 => x"f0050c80",
  9045 => x"0b8c08f4",
  9046 => x"050c8c08",
  9047 => x"8c05088c",
  9048 => x"08900508",
  9049 => x"5654738c",
  9050 => x"08f0050c",
  9051 => x"748c08f4",
  9052 => x"050c8c08",
  9053 => x"f8058c08",
  9054 => x"f0055656",
  9055 => x"88705475",
  9056 => x"53765254",
  9057 => x"fdf7883f",
  9058 => x"a00b8c08",
  9059 => x"94050831",
  9060 => x"8c08ec05",
  9061 => x"0c8c08ec",
  9062 => x"05088024",
  9063 => x"9d38800b",
  9064 => x"8c08f005",
  9065 => x"0c8c08ec",
  9066 => x"0508308c",
  9067 => x"08f80508",
  9068 => x"712a8c08",
  9069 => x"f4050c54",
  9070 => x"b9398c08",
  9071 => x"f805088c",
  9072 => x"08ec0508",
  9073 => x"2b8c08e8",
  9074 => x"050c8c08",
  9075 => x"f805088c",
  9076 => x"08940508",
  9077 => x"2a8c08f0",
  9078 => x"050c8c08",
  9079 => x"fc05088c",
  9080 => x"08940508",
  9081 => x"2a708c08",
  9082 => x"e8050807",
  9083 => x"8c08f405",
  9084 => x"0c548c08",
  9085 => x"f005088c",
  9086 => x"08f40508",
  9087 => x"8c088805",
  9088 => x"08585654",
  9089 => x"73760c74",
  9090 => x"84170c8c",
  9091 => x"08880508",
  9092 => x"800c8d3d",
  9093 => x"0d8c0c04",
  9094 => x"8c08028c",
  9095 => x"0cc73d0d",
  9096 => x"8c088c05",
  9097 => x"08559015",
  9098 => x"088c1608",
  9099 => x"5656748c",
  9100 => x"08f0050c",
  9101 => x"758c08f4",
  9102 => x"050c8c08",
  9103 => x"8c050884",
  9104 => x"11088c08",
  9105 => x"ec050c55",
  9106 => x"800b8c08",
  9107 => x"e8050c8c",
  9108 => x"088c0508",
  9109 => x"518fb83f",
  9110 => x"80085574",
  9111 => x"802eaa38",
  9112 => x"8fff0b8c",
  9113 => x"08e8050c",
  9114 => x"8c08f005",
  9115 => x"08a08080",
  9116 => x"078c08f4",
  9117 => x"05088007",
  9118 => x"5755748c",
  9119 => x"08f0050c",
  9120 => x"758c08f4",
  9121 => x"050c8d80",
  9122 => x"398c088c",
  9123 => x"0508518e",
  9124 => x"ca3f8008",
  9125 => x"5574802e",
  9126 => x"9c388fff",
  9127 => x"0b8c08e8",
  9128 => x"050c8055",
  9129 => x"8056748c",
  9130 => x"08f0050c",
  9131 => x"758c08f4",
  9132 => x"050c8cd4",
  9133 => x"398c088c",
  9134 => x"0508518d",
  9135 => x"ea3f8008",
  9136 => x"5574802e",
  9137 => x"9b38800b",
  9138 => x"8c08e805",
  9139 => x"0c805580",
  9140 => x"56748c08",
  9141 => x"f0050c75",
  9142 => x"8c08f405",
  9143 => x"0c8ca939",
  9144 => x"8c08f005",
  9145 => x"08708c08",
  9146 => x"f4050807",
  9147 => x"5155748b",
  9148 => x"38800b8c",
  9149 => x"08e8050c",
  9150 => x"8c8e398c",
  9151 => x"088c0508",
  9152 => x"55881508",
  9153 => x"f8822586",
  9154 => x"fc388c08",
  9155 => x"8c0508f8",
  9156 => x"820b8812",
  9157 => x"08318c08",
  9158 => x"e4050c55",
  9159 => x"800b8c08",
  9160 => x"e8050cb8",
  9161 => x"0b8c08e4",
  9162 => x"05082594",
  9163 => x"38805580",
  9164 => x"56748c08",
  9165 => x"f0050c75",
  9166 => x"8c08f405",
  9167 => x"0c82a339",
  9168 => x"800b8c08",
  9169 => x"e0050c8c",
  9170 => x"08d80557",
  9171 => x"8055810b",
  9172 => x"8c08e405",
  9173 => x"08555674",
  9174 => x"52755376",
  9175 => x"51fded89",
  9176 => x"3f8c08d8",
  9177 => x"05088c08",
  9178 => x"dc050857",
  9179 => x"55748c08",
  9180 => x"d0050c75",
  9181 => x"8c08d405",
  9182 => x"0cff56ff",
  9183 => x"57758c08",
  9184 => x"c8050c76",
  9185 => x"8c08cc05",
  9186 => x"0c8c08d4",
  9187 => x"05088c08",
  9188 => x"cc050870",
  9189 => x"12708c08",
  9190 => x"c4050c52",
  9191 => x"5657810b",
  9192 => x"8c08ffbc",
  9193 => x"050c8c08",
  9194 => x"c405088c",
  9195 => x"08d40508",
  9196 => x"58567676",
  9197 => x"26893880",
  9198 => x"0b8c08ff",
  9199 => x"bc050c8c",
  9200 => x"08d00508",
  9201 => x"8c08c805",
  9202 => x"08701270",
  9203 => x"8c08c005",
  9204 => x"0c8c08c0",
  9205 => x"05088c08",
  9206 => x"ffbc0508",
  9207 => x"11708c08",
  9208 => x"c0050c8c",
  9209 => x"08c00508",
  9210 => x"708c08f0",
  9211 => x"0508068c",
  9212 => x"08c40508",
  9213 => x"708c08f4",
  9214 => x"05080672",
  9215 => x"70720751",
  9216 => x"52575252",
  9217 => x"52525a52",
  9218 => x"57557680",
  9219 => x"2e883881",
  9220 => x"0b8c08e0",
  9221 => x"050c8c08",
  9222 => x"d8058c08",
  9223 => x"e4050855",
  9224 => x"578c08f0",
  9225 => x"05088c08",
  9226 => x"f4050857",
  9227 => x"55745275",
  9228 => x"537651f9",
  9229 => x"ec3f8c08",
  9230 => x"d805088c",
  9231 => x"08dc0508",
  9232 => x"8c08e005",
  9233 => x"089f2c8c",
  9234 => x"08e00508",
  9235 => x"71707507",
  9236 => x"8c08f005",
  9237 => x"0c737207",
  9238 => x"8c08f405",
  9239 => x"0c59595b",
  9240 => x"59578c08",
  9241 => x"f0050880",
  9242 => x"06708c08",
  9243 => x"ffb4050c",
  9244 => x"8c08f405",
  9245 => x"0881ff06",
  9246 => x"708c08ff",
  9247 => x"b8050c57",
  9248 => x"558c08ff",
  9249 => x"b405088c",
  9250 => x"08ffb805",
  9251 => x"08575574",
  9252 => x"8c08ffb4",
  9253 => x"050c758c",
  9254 => x"08ffb805",
  9255 => x"0c8c08ff",
  9256 => x"b4050856",
  9257 => x"7581eb38",
  9258 => x"8c08ffb8",
  9259 => x"05085776",
  9260 => x"81802e09",
  9261 => x"810681da",
  9262 => x"388c08f0",
  9263 => x"0508982b",
  9264 => x"8c08f405",
  9265 => x"08882a70",
  9266 => x"72078c08",
  9267 => x"f0050888",
  9268 => x"2a718106",
  9269 => x"51585858",
  9270 => x"5874802e",
  9271 => x"82e4388c",
  9272 => x"08f00508",
  9273 => x"8c08f405",
  9274 => x"08575574",
  9275 => x"8c08ffac",
  9276 => x"050c758c",
  9277 => x"08ffb005",
  9278 => x"0c805681",
  9279 => x"8057758c",
  9280 => x"08ffa405",
  9281 => x"0c768c08",
  9282 => x"ffa8050c",
  9283 => x"8c08ffb0",
  9284 => x"05088c08",
  9285 => x"ffa80508",
  9286 => x"7012708c",
  9287 => x"08ffa005",
  9288 => x"0c525657",
  9289 => x"810b8c08",
  9290 => x"ff98050c",
  9291 => x"8c08ffa0",
  9292 => x"05088c08",
  9293 => x"ffb00508",
  9294 => x"58567676",
  9295 => x"26893880",
  9296 => x"0b8c08ff",
  9297 => x"98050c8c",
  9298 => x"08ffac05",
  9299 => x"088c08ff",
  9300 => x"a4050870",
  9301 => x"12708c08",
  9302 => x"ff9c050c",
  9303 => x"8c08ff9c",
  9304 => x"05088c08",
  9305 => x"ff980508",
  9306 => x"11708c08",
  9307 => x"ff9c050c",
  9308 => x"525a5257",
  9309 => x"558c08ff",
  9310 => x"9c05088c",
  9311 => x"08ffa005",
  9312 => x"08575574",
  9313 => x"8c08f005",
  9314 => x"0c758c08",
  9315 => x"f4050c81",
  9316 => x"b1398c08",
  9317 => x"f005088c",
  9318 => x"08f40508",
  9319 => x"5856758c",
  9320 => x"08ff9005",
  9321 => x"0c768c08",
  9322 => x"ff94050c",
  9323 => x"805580ff",
  9324 => x"56748c08",
  9325 => x"ff88050c",
  9326 => x"758c08ff",
  9327 => x"8c050c8c",
  9328 => x"08ff9405",
  9329 => x"088c08ff",
  9330 => x"8c050870",
  9331 => x"12708c08",
  9332 => x"ff84050c",
  9333 => x"52585681",
  9334 => x"0b8c08fe",
  9335 => x"fc050c8c",
  9336 => x"08ff8405",
  9337 => x"088c08ff",
  9338 => x"94050857",
  9339 => x"55757526",
  9340 => x"8938800b",
  9341 => x"8c08fefc",
  9342 => x"050c8c08",
  9343 => x"ff900508",
  9344 => x"8c08ff88",
  9345 => x"05087012",
  9346 => x"708c08ff",
  9347 => x"80050c8c",
  9348 => x"08ff8005",
  9349 => x"088c08fe",
  9350 => x"fc050811",
  9351 => x"708c08ff",
  9352 => x"80050c53",
  9353 => x"59525657",
  9354 => x"8c08ff80",
  9355 => x"05088c08",
  9356 => x"ff840508",
  9357 => x"5755748c",
  9358 => x"08f0050c",
  9359 => x"758c08f4",
  9360 => x"050c8c08",
  9361 => x"f00508f0",
  9362 => x"0a268338",
  9363 => x"8d398c08",
  9364 => x"e8050881",
  9365 => x"058c08e8",
  9366 => x"050c8c08",
  9367 => x"f0050898",
  9368 => x"2b8c08f4",
  9369 => x"0508882a",
  9370 => x"7072078c",
  9371 => x"08f00508",
  9372 => x"882a5858",
  9373 => x"5858748c",
  9374 => x"08f0050c",
  9375 => x"758c08f4",
  9376 => x"050c8584",
  9377 => x"398c088c",
  9378 => x"05085587",
  9379 => x"ff0b8816",
  9380 => x"08259c38",
  9381 => x"8fff0b8c",
  9382 => x"08e8050c",
  9383 => x"80558056",
  9384 => x"748c08f0",
  9385 => x"050c758c",
  9386 => x"08f4050c",
  9387 => x"84da398c",
  9388 => x"088c0508",
  9389 => x"88110887",
  9390 => x"ff058c08",
  9391 => x"e8050c8c",
  9392 => x"08f00508",
  9393 => x"8006708c",
  9394 => x"08fef405",
  9395 => x"0c8c08f4",
  9396 => x"050881ff",
  9397 => x"06708c08",
  9398 => x"fef8050c",
  9399 => x"5957558c",
  9400 => x"08fef405",
  9401 => x"088c08fe",
  9402 => x"f8050857",
  9403 => x"55748c08",
  9404 => x"fef4050c",
  9405 => x"758c08fe",
  9406 => x"f8050c8c",
  9407 => x"08fef405",
  9408 => x"08567581",
  9409 => x"eb388c08",
  9410 => x"fef80508",
  9411 => x"57768180",
  9412 => x"2e098106",
  9413 => x"81da388c",
  9414 => x"08f00508",
  9415 => x"982b8c08",
  9416 => x"f4050888",
  9417 => x"2a707207",
  9418 => x"8c08f005",
  9419 => x"08882a71",
  9420 => x"81065158",
  9421 => x"58585874",
  9422 => x"802e82e4",
  9423 => x"388c08f0",
  9424 => x"05088c08",
  9425 => x"f4050857",
  9426 => x"55748c08",
  9427 => x"feec050c",
  9428 => x"758c08fe",
  9429 => x"f0050c80",
  9430 => x"56818057",
  9431 => x"758c08fe",
  9432 => x"e4050c76",
  9433 => x"8c08fee8",
  9434 => x"050c8c08",
  9435 => x"fef00508",
  9436 => x"8c08fee8",
  9437 => x"05087012",
  9438 => x"708c08fe",
  9439 => x"e0050c52",
  9440 => x"5657810b",
  9441 => x"8c08fed8",
  9442 => x"050c8c08",
  9443 => x"fee00508",
  9444 => x"8c08fef0",
  9445 => x"05085856",
  9446 => x"76762689",
  9447 => x"38800b8c",
  9448 => x"08fed805",
  9449 => x"0c8c08fe",
  9450 => x"ec05088c",
  9451 => x"08fee405",
  9452 => x"08701270",
  9453 => x"8c08fedc",
  9454 => x"050c8c08",
  9455 => x"fedc0508",
  9456 => x"8c08fed8",
  9457 => x"05081170",
  9458 => x"8c08fedc",
  9459 => x"050c525a",
  9460 => x"5257558c",
  9461 => x"08fedc05",
  9462 => x"088c08fe",
  9463 => x"e0050857",
  9464 => x"55748c08",
  9465 => x"f0050c75",
  9466 => x"8c08f405",
  9467 => x"0c81b139",
  9468 => x"8c08f005",
  9469 => x"088c08f4",
  9470 => x"05085856",
  9471 => x"758c08fe",
  9472 => x"d0050c76",
  9473 => x"8c08fed4",
  9474 => x"050c8055",
  9475 => x"80ff5674",
  9476 => x"8c08fec8",
  9477 => x"050c758c",
  9478 => x"08fecc05",
  9479 => x"0c8c08fe",
  9480 => x"d405088c",
  9481 => x"08fecc05",
  9482 => x"08701270",
  9483 => x"8c08fec4",
  9484 => x"050c5258",
  9485 => x"56810b8c",
  9486 => x"08febc05",
  9487 => x"0c8c08fe",
  9488 => x"c405088c",
  9489 => x"08fed405",
  9490 => x"08575575",
  9491 => x"75268938",
  9492 => x"800b8c08",
  9493 => x"febc050c",
  9494 => x"8c08fed0",
  9495 => x"05088c08",
  9496 => x"fec80508",
  9497 => x"7012708c",
  9498 => x"08fec005",
  9499 => x"0c8c08fe",
  9500 => x"c005088c",
  9501 => x"08febc05",
  9502 => x"0811708c",
  9503 => x"08fec005",
  9504 => x"0c535952",
  9505 => x"56578c08",
  9506 => x"fec00508",
  9507 => x"8c08fec4",
  9508 => x"05085755",
  9509 => x"748c08f0",
  9510 => x"050c758c",
  9511 => x"08f4050c",
  9512 => x"8c08f005",
  9513 => x"08f80a26",
  9514 => x"8338b539",
  9515 => x"8c08f005",
  9516 => x"089f2b8c",
  9517 => x"08f40508",
  9518 => x"812a7072",
  9519 => x"078c08f0",
  9520 => x"0508812a",
  9521 => x"58585858",
  9522 => x"748c08f0",
  9523 => x"050c758c",
  9524 => x"08f4050c",
  9525 => x"8c08e805",
  9526 => x"0881058c",
  9527 => x"08e8050c",
  9528 => x"8c08f005",
  9529 => x"08982b8c",
  9530 => x"08f40508",
  9531 => x"882a7072",
  9532 => x"078c08f0",
  9533 => x"0508882a",
  9534 => x"58585858",
  9535 => x"748c08f0",
  9536 => x"050c758c",
  9537 => x"08f4050c",
  9538 => x"8c08f005",
  9539 => x"08bfffff",
  9540 => x"068c08f8",
  9541 => x"050c8c08",
  9542 => x"f40508ff",
  9543 => x"068c08fc",
  9544 => x"050c8c08",
  9545 => x"e8050856",
  9546 => x"80708006",
  9547 => x"778fff06",
  9548 => x"70942b53",
  9549 => x"5a585580",
  9550 => x"0b8c08f8",
  9551 => x"05087607",
  9552 => x"8c08f805",
  9553 => x"0c708c08",
  9554 => x"fc050807",
  9555 => x"8c08fc05",
  9556 => x"0c8c08ec",
  9557 => x"05085156",
  9558 => x"80708006",
  9559 => x"77810670",
  9560 => x"9f2b535a",
  9561 => x"5855800b",
  9562 => x"8c08f805",
  9563 => x"0876078c",
  9564 => x"08f8050c",
  9565 => x"708c08fc",
  9566 => x"0508078c",
  9567 => x"08fc050c",
  9568 => x"568c08f8",
  9569 => x"05088c08",
  9570 => x"fc05088c",
  9571 => x"08880508",
  9572 => x"59575574",
  9573 => x"770c7584",
  9574 => x"180c8c08",
  9575 => x"88050880",
  9576 => x"0cbb3d0d",
  9577 => x"8c0c048c",
  9578 => x"08028c0c",
  9579 => x"ff3d0d80",
  9580 => x"0b8c08fc",
  9581 => x"050c8c08",
  9582 => x"88050851",
  9583 => x"7008822e",
  9584 => x"09810688",
  9585 => x"38810b8c",
  9586 => x"08fc050c",
  9587 => x"8c08fc05",
  9588 => x"0870800c",
  9589 => x"51833d0d",
  9590 => x"8c0c048c",
  9591 => x"08028c0c",
  9592 => x"ff3d0d80",
  9593 => x"0b8c08fc",
  9594 => x"050c8c08",
  9595 => x"88050851",
  9596 => x"7008842e",
  9597 => x"09810688",
  9598 => x"38810b8c",
  9599 => x"08fc050c",
  9600 => x"8c08fc05",
  9601 => x"0870800c",
  9602 => x"51833d0d",
  9603 => x"8c0c048c",
  9604 => x"08028c0c",
  9605 => x"ff3d0d80",
  9606 => x"0b8c08fc",
  9607 => x"050c8c08",
  9608 => x"88050851",
  9609 => x"7008802e",
  9610 => x"8f388c08",
  9611 => x"88050851",
  9612 => x"7008812e",
  9613 => x"83388839",
  9614 => x"810b8c08",
  9615 => x"fc050c8c",
  9616 => x"08fc0508",
  9617 => x"70800c51",
  9618 => x"833d0d8c",
  9619 => x"0c048c08",
  9620 => x"028c0cf8",
  9621 => x"3d0d8c08",
  9622 => x"88050870",
  9623 => x"08bfffff",
  9624 => x"068c08f8",
  9625 => x"050c8411",
  9626 => x"08ff068c",
  9627 => x"08fc050c",
  9628 => x"8c088805",
  9629 => x"08700894",
  9630 => x"2a545451",
  9631 => x"80728fff",
  9632 => x"068c08f4",
  9633 => x"050c8c08",
  9634 => x"88050870",
  9635 => x"089f2a54",
  9636 => x"54518072",
  9637 => x"81068c08",
  9638 => x"f0050c8c",
  9639 => x"088c0508",
  9640 => x"8c08f005",
  9641 => x"0884120c",
  9642 => x"51518c08",
  9643 => x"f4050881",
  9644 => x"bd388c08",
  9645 => x"f8050870",
  9646 => x"8c08fc05",
  9647 => x"08075151",
  9648 => x"708d388c",
  9649 => x"088c0508",
  9650 => x"5182710c",
  9651 => x"82d8398c",
  9652 => x"088c0508",
  9653 => x"8c08f405",
  9654 => x"08f88205",
  9655 => x"88120c8c",
  9656 => x"08fc0508",
  9657 => x"982a8c08",
  9658 => x"f8050888",
  9659 => x"2b707207",
  9660 => x"8c08fc05",
  9661 => x"08882b56",
  9662 => x"53555551",
  9663 => x"708c08f8",
  9664 => x"050c718c",
  9665 => x"08fc050c",
  9666 => x"8c088c05",
  9667 => x"08518371",
  9668 => x"0c8c08f8",
  9669 => x"0508f00a",
  9670 => x"26b7388c",
  9671 => x"08fc0508",
  9672 => x"9f2a8c08",
  9673 => x"f8050810",
  9674 => x"7072078c",
  9675 => x"08fc0508",
  9676 => x"10555354",
  9677 => x"54708c08",
  9678 => x"f8050c71",
  9679 => x"8c08fc05",
  9680 => x"0c8c088c",
  9681 => x"05088811",
  9682 => x"08ff0588",
  9683 => x"120c51c1",
  9684 => x"398c088c",
  9685 => x"0508538c",
  9686 => x"08f80508",
  9687 => x"8c08fc05",
  9688 => x"08535170",
  9689 => x"8c140c71",
  9690 => x"90140c81",
  9691 => x"b9398c08",
  9692 => x"f405088f",
  9693 => x"ff2e0981",
  9694 => x"0680e238",
  9695 => x"8c08f805",
  9696 => x"08708c08",
  9697 => x"fc050807",
  9698 => x"5151708d",
  9699 => x"388c088c",
  9700 => x"05085184",
  9701 => x"710c818e",
  9702 => x"398c08f8",
  9703 => x"0508932a",
  9704 => x"52807281",
  9705 => x"06515170",
  9706 => x"802e8c38",
  9707 => x"8c088c05",
  9708 => x"08518171",
  9709 => x"0c8a398c",
  9710 => x"088c0508",
  9711 => x"5180710c",
  9712 => x"8c088c05",
  9713 => x"08538c08",
  9714 => x"f805088c",
  9715 => x"08fc0508",
  9716 => x"5351708c",
  9717 => x"140c7190",
  9718 => x"140c80ca",
  9719 => x"398c088c",
  9720 => x"05088c08",
  9721 => x"f40508f8",
  9722 => x"81058812",
  9723 => x"0c8c088c",
  9724 => x"05085151",
  9725 => x"83710c8c",
  9726 => x"088c0508",
  9727 => x"8c08fc05",
  9728 => x"08982a8c",
  9729 => x"08f80508",
  9730 => x"882b7072",
  9731 => x"078c08fc",
  9732 => x"0508882b",
  9733 => x"71880a07",
  9734 => x"8c160c70",
  9735 => x"80079016",
  9736 => x"0c565455",
  9737 => x"55558a3d",
  9738 => x"0d8c0c04",
  9739 => x"8c08028c",
  9740 => x"0cf03d0d",
  9741 => x"8c088805",
  9742 => x"085187b7",
  9743 => x"3f800852",
  9744 => x"7192388c",
  9745 => x"088c0508",
  9746 => x"5187a83f",
  9747 => x"80085271",
  9748 => x"83388b39",
  9749 => x"810b8c08",
  9750 => x"fc050c86",
  9751 => x"a1398c08",
  9752 => x"88050851",
  9753 => x"86d93f80",
  9754 => x"08527180",
  9755 => x"2eaf388c",
  9756 => x"088c0508",
  9757 => x"5186c83f",
  9758 => x"80085271",
  9759 => x"802e9e38",
  9760 => x"8c088c05",
  9761 => x"088c0888",
  9762 => x"05088412",
  9763 => x"08841208",
  9764 => x"31708c08",
  9765 => x"fc050c52",
  9766 => x"545285e2",
  9767 => x"398c0888",
  9768 => x"05085186",
  9769 => x"9a3f8008",
  9770 => x"5271802e",
  9771 => x"ab388c08",
  9772 => x"88050852",
  9773 => x"84120880",
  9774 => x"2e8a38ff",
  9775 => x"0b8c08f8",
  9776 => x"050c8839",
  9777 => x"810b8c08",
  9778 => x"f8050c8c",
  9779 => x"08f80508",
  9780 => x"8c08fc05",
  9781 => x"0c85a739",
  9782 => x"8c088c05",
  9783 => x"085185df",
  9784 => x"3f800852",
  9785 => x"71802eab",
  9786 => x"388c088c",
  9787 => x"05085284",
  9788 => x"1208802e",
  9789 => x"8a38810b",
  9790 => x"8c08f405",
  9791 => x"0c8839ff",
  9792 => x"0b8c08f4",
  9793 => x"050c8c08",
  9794 => x"f405088c",
  9795 => x"08fc050c",
  9796 => x"84ec398c",
  9797 => x"08880508",
  9798 => x"5184f03f",
  9799 => x"80085271",
  9800 => x"802e9c38",
  9801 => x"8c088c05",
  9802 => x"085184df",
  9803 => x"3f800852",
  9804 => x"71802e8b",
  9805 => x"38800b8c",
  9806 => x"08fc050c",
  9807 => x"84c0398c",
  9808 => x"08880508",
  9809 => x"5184c43f",
  9810 => x"80085271",
  9811 => x"802eab38",
  9812 => x"8c088c05",
  9813 => x"08528412",
  9814 => x"08802e8a",
  9815 => x"38810b8c",
  9816 => x"08f0050c",
  9817 => x"8839ff0b",
  9818 => x"8c08f005",
  9819 => x"0c8c08f0",
  9820 => x"05088c08",
  9821 => x"fc050c84",
  9822 => x"85398c08",
  9823 => x"8c050851",
  9824 => x"84893f80",
  9825 => x"08527180",
  9826 => x"2eab388c",
  9827 => x"08880508",
  9828 => x"52841208",
  9829 => x"802e8a38",
  9830 => x"ff0b8c08",
  9831 => x"ec050c88",
  9832 => x"39810b8c",
  9833 => x"08ec050c",
  9834 => x"8c08ec05",
  9835 => x"088c08fc",
  9836 => x"050c83ca",
  9837 => x"398c0888",
  9838 => x"05088c08",
  9839 => x"8c050853",
  9840 => x"53841308",
  9841 => x"8413082e",
  9842 => x"ab388c08",
  9843 => x"88050852",
  9844 => x"84120880",
  9845 => x"2e8a38ff",
  9846 => x"0b8c08e8",
  9847 => x"050c8839",
  9848 => x"810b8c08",
  9849 => x"e8050c8c",
  9850 => x"08e80508",
  9851 => x"8c08fc05",
  9852 => x"0c838b39",
  9853 => x"8c088805",
  9854 => x"088c088c",
  9855 => x"05085353",
  9856 => x"88120888",
  9857 => x"140825ab",
  9858 => x"388c0888",
  9859 => x"05085284",
  9860 => x"1208802e",
  9861 => x"8a38ff0b",
  9862 => x"8c08e405",
  9863 => x"0c883981",
  9864 => x"0b8c08e4",
  9865 => x"050c8c08",
  9866 => x"e405088c",
  9867 => x"08fc050c",
  9868 => x"82cc398c",
  9869 => x"08880508",
  9870 => x"8c088c05",
  9871 => x"08535388",
  9872 => x"13088813",
  9873 => x"0825ab38",
  9874 => x"8c088805",
  9875 => x"08528412",
  9876 => x"08802e8a",
  9877 => x"38810b8c",
  9878 => x"08e0050c",
  9879 => x"8839ff0b",
  9880 => x"8c08e005",
  9881 => x"0c8c08e0",
  9882 => x"05088c08",
  9883 => x"fc050c82",
  9884 => x"8d398c08",
  9885 => x"8805088c",
  9886 => x"08dc050c",
  9887 => x"8c088c05",
  9888 => x"088c08d8",
  9889 => x"050c8c08",
  9890 => x"dc05088c",
  9891 => x"08d80508",
  9892 => x"54528c12",
  9893 => x"088c1408",
  9894 => x"26b1388c",
  9895 => x"08dc0508",
  9896 => x"8c08d805",
  9897 => x"0854528c",
  9898 => x"12088c14",
  9899 => x"082e0981",
  9900 => x"0680c238",
  9901 => x"8c08dc05",
  9902 => x"088c08d8",
  9903 => x"05085452",
  9904 => x"90120890",
  9905 => x"14082683",
  9906 => x"38ab398c",
  9907 => x"08880508",
  9908 => x"52841208",
  9909 => x"802e8a38",
  9910 => x"ff0b8c08",
  9911 => x"d4050c88",
  9912 => x"39810b8c",
  9913 => x"08d4050c",
  9914 => x"8c08d405",
  9915 => x"088c08fc",
  9916 => x"050c818a",
  9917 => x"398c088c",
  9918 => x"05088c08",
  9919 => x"d0050c8c",
  9920 => x"08880508",
  9921 => x"8c08cc05",
  9922 => x"0c8c08d0",
  9923 => x"05088c08",
  9924 => x"cc050854",
  9925 => x"528c1208",
  9926 => x"8c140826",
  9927 => x"b1388c08",
  9928 => x"d005088c",
  9929 => x"08cc0508",
  9930 => x"54528c12",
  9931 => x"088c1408",
  9932 => x"2e098106",
  9933 => x"80c1388c",
  9934 => x"08d00508",
  9935 => x"8c08cc05",
  9936 => x"08545290",
  9937 => x"12089014",
  9938 => x"08268338",
  9939 => x"aa398c08",
  9940 => x"88050852",
  9941 => x"84120880",
  9942 => x"2e8a3881",
  9943 => x"0b8c08c8",
  9944 => x"050c8839",
  9945 => x"ff0b8c08",
  9946 => x"c8050c8c",
  9947 => x"08c80508",
  9948 => x"8c08fc05",
  9949 => x"0c883980",
  9950 => x"0b8c08fc",
  9951 => x"050c8c08",
  9952 => x"fc050880",
  9953 => x"0c923d0d",
  9954 => x"8c0c048c",
  9955 => x"08028c0c",
  9956 => x"ff3d0d80",
  9957 => x"0b8c08fc",
  9958 => x"050c8c08",
  9959 => x"88050851",
  9960 => x"7008822e",
  9961 => x"09810688",
  9962 => x"38810b8c",
  9963 => x"08fc050c",
  9964 => x"8c08fc05",
  9965 => x"0870800c",
  9966 => x"51833d0d",
  9967 => x"8c0c048c",
  9968 => x"08028c0c",
  9969 => x"ff3d0d80",
  9970 => x"0b8c08fc",
  9971 => x"050c8c08",
  9972 => x"88050851",
  9973 => x"7008842e",
  9974 => x"09810688",
  9975 => x"38810b8c",
  9976 => x"08fc050c",
  9977 => x"8c08fc05",
  9978 => x"0870800c",
  9979 => x"51833d0d",
  9980 => x"8c0c048c",
  9981 => x"08028c0c",
  9982 => x"ff3d0d80",
  9983 => x"0b8c08fc",
  9984 => x"050c8c08",
  9985 => x"88050851",
  9986 => x"7008802e",
  9987 => x"8f388c08",
  9988 => x"88050851",
  9989 => x"7008812e",
  9990 => x"83388839",
  9991 => x"810b8c08",
  9992 => x"fc050c8c",
  9993 => x"08fc0508",
  9994 => x"70800c51",
  9995 => x"833d0d8c",
  9996 => x"0c04ff3d",
  9997 => x"0d82d0ac",
  9998 => x"0bfc0570",
  9999 => x"08525270",
 10000 => x"ff2e9138",
 10001 => x"702dfc12",
 10002 => x"70085252",
 10003 => x"70ff2e09",
 10004 => x"8106f138",
 10005 => x"833d0d04",
 10006 => x"04fdd084",
 10007 => x"3f040000",
 10008 => x"48656c6c",
 10009 => x"6f20776f",
 10010 => x"726c6421",
 10011 => x"3a202563",
 10012 => x"0a000000",
 10013 => x"00000040",
 10014 => x"20202020",
 10015 => x"20202020",
 10016 => x"20202020",
 10017 => x"20202020",
 10018 => x"30303030",
 10019 => x"30303030",
 10020 => x"30303030",
 10021 => x"30303030",
 10022 => x"000013a9",
 10023 => x"00000f58",
 10024 => x"00000f58",
 10025 => x"0000139f",
 10026 => x"00000f58",
 10027 => x"00000f58",
 10028 => x"00000f58",
 10029 => x"00000f58",
 10030 => x"00000f58",
 10031 => x"00000f58",
 10032 => x"00000f2f",
 10033 => x"0000133e",
 10034 => x"00000f58",
 10035 => x"00000f41",
 10036 => x"000010e1",
 10037 => x"00000f58",
 10038 => x"0000136c",
 10039 => x"0000134a",
 10040 => x"0000134a",
 10041 => x"0000134a",
 10042 => x"0000134a",
 10043 => x"0000134a",
 10044 => x"0000134a",
 10045 => x"0000134a",
 10046 => x"0000134a",
 10047 => x"0000134a",
 10048 => x"00000f58",
 10049 => x"00000f58",
 10050 => x"00000f58",
 10051 => x"00000f58",
 10052 => x"00000f58",
 10053 => x"00000f58",
 10054 => x"00000f58",
 10055 => x"00000f58",
 10056 => x"00000f58",
 10057 => x"00001231",
 10058 => x"00000ef7",
 10059 => x"000011ba",
 10060 => x"00000f58",
 10061 => x"000011ba",
 10062 => x"00000f58",
 10063 => x"00000f58",
 10064 => x"00000f58",
 10065 => x"00000f58",
 10066 => x"00001377",
 10067 => x"00000f58",
 10068 => x"00000f58",
 10069 => x"00000ec4",
 10070 => x"00000f58",
 10071 => x"00000f58",
 10072 => x"00000f58",
 10073 => x"000012c2",
 10074 => x"00000f58",
 10075 => x"00000c12",
 10076 => x"00000f58",
 10077 => x"00000f58",
 10078 => x"0000127b",
 10079 => x"00000f58",
 10080 => x"00000f58",
 10081 => x"00000f58",
 10082 => x"00000f58",
 10083 => x"00000f58",
 10084 => x"00000f58",
 10085 => x"00000f58",
 10086 => x"00000f58",
 10087 => x"00000f58",
 10088 => x"00000f58",
 10089 => x"00001231",
 10090 => x"00000efb",
 10091 => x"000011ba",
 10092 => x"000011ba",
 10093 => x"000011ba",
 10094 => x"000011af",
 10095 => x"00000efb",
 10096 => x"00000f58",
 10097 => x"00000f58",
 10098 => x"000010c3",
 10099 => x"00000f58",
 10100 => x"00001313",
 10101 => x"00000ec8",
 10102 => x"00001124",
 10103 => x"00000f4e",
 10104 => x"00000f58",
 10105 => x"000012c2",
 10106 => x"00000f58",
 10107 => x"00000c16",
 10108 => x"00000f58",
 10109 => x"00000f58",
 10110 => x"00001381",
 10111 => x"62756720",
 10112 => x"696e2076",
 10113 => x"66707269",
 10114 => x"6e74663a",
 10115 => x"20626164",
 10116 => x"20626173",
 10117 => x"65000000",
 10118 => x"30313233",
 10119 => x"34353637",
 10120 => x"38396162",
 10121 => x"63646566",
 10122 => x"00000000",
 10123 => x"496e6600",
 10124 => x"30313233",
 10125 => x"34353637",
 10126 => x"38394142",
 10127 => x"43444546",
 10128 => x"00000000",
 10129 => x"30000000",
 10130 => x"2e000000",
 10131 => x"4e614e00",
 10132 => x"286e756c",
 10133 => x"6c290000",
 10134 => x"432d5554",
 10135 => x"462d3800",
 10136 => x"432d534a",
 10137 => x"49530000",
 10138 => x"432d4555",
 10139 => x"434a5000",
 10140 => x"432d4a49",
 10141 => x"53000000",
 10142 => x"496e6669",
 10143 => x"6e697479",
 10144 => x"00000000",
 10145 => x"00002fbc",
 10146 => x"00002fbc",
 10147 => x"00002fa6",
 10148 => x"00002abb",
 10149 => x"00002fab",
 10150 => x"00002ac0",
 10151 => x"43000000",
 10152 => x"49534f2d",
 10153 => x"38383539",
 10154 => x"2d310000",
 10155 => x"00009e48",
 10156 => x"00009e40",
 10157 => x"00009e40",
 10158 => x"00009e40",
 10159 => x"00009e40",
 10160 => x"00009e40",
 10161 => x"00009e40",
 10162 => x"00009e40",
 10163 => x"00009e40",
 10164 => x"00009e40",
 10165 => x"ffffffff",
 10166 => x"ffffffff",
 10167 => x"3c9cd2b2",
 10168 => x"97d889bc",
 10169 => x"3949f623",
 10170 => x"d5a8a733",
 10171 => x"32a50ffd",
 10172 => x"44f4a73d",
 10173 => x"255bba08",
 10174 => x"cf8c979d",
 10175 => x"0ac80628",
 10176 => x"64ac6f43",
 10177 => x"4341c379",
 10178 => x"37e08000",
 10179 => x"4693b8b5",
 10180 => x"b5056e17",
 10181 => x"4d384f03",
 10182 => x"e93ff9f5",
 10183 => x"5a827748",
 10184 => x"f9301d32",
 10185 => x"75154fdd",
 10186 => x"7f73bf3c",
 10187 => x"3ff00000",
 10188 => x"00000000",
 10189 => x"40240000",
 10190 => x"00000000",
 10191 => x"40590000",
 10192 => x"00000000",
 10193 => x"408f4000",
 10194 => x"00000000",
 10195 => x"40c38800",
 10196 => x"00000000",
 10197 => x"40f86a00",
 10198 => x"00000000",
 10199 => x"412e8480",
 10200 => x"00000000",
 10201 => x"416312d0",
 10202 => x"00000000",
 10203 => x"4197d784",
 10204 => x"00000000",
 10205 => x"41cdcd65",
 10206 => x"00000000",
 10207 => x"4202a05f",
 10208 => x"20000000",
 10209 => x"42374876",
 10210 => x"e8000000",
 10211 => x"426d1a94",
 10212 => x"a2000000",
 10213 => x"42a2309c",
 10214 => x"e5400000",
 10215 => x"42d6bcc4",
 10216 => x"1e900000",
 10217 => x"430c6bf5",
 10218 => x"26340000",
 10219 => x"4341c379",
 10220 => x"37e08000",
 10221 => x"43763457",
 10222 => x"85d8a000",
 10223 => x"43abc16d",
 10224 => x"674ec800",
 10225 => x"43e158e4",
 10226 => x"60913d00",
 10227 => x"4415af1d",
 10228 => x"78b58c40",
 10229 => x"444b1ae4",
 10230 => x"d6e2ef50",
 10231 => x"4480f0cf",
 10232 => x"064dd592",
 10233 => x"44b52d02",
 10234 => x"c7e14af6",
 10235 => x"44ea7843",
 10236 => x"79d99db4",
 10237 => x"00000005",
 10238 => x"00000019",
 10239 => x"0000007d",
 10240 => x"64756d6d",
 10241 => x"792e6578",
 10242 => x"65000000",
 10243 => x"00000000",
 10244 => x"00000000",
 10245 => x"00000000",
 10246 => x"00000000",
 10247 => x"00000000",
 10248 => x"00ffffff",
 10249 => x"ff00ffff",
 10250 => x"ffff00ff",
 10251 => x"ffffff00",
 10252 => x"00000000",
 10253 => x"00000000",
 10254 => x"00000000",
 10255 => x"0000a834",
 10256 => x"0000a044",
 10257 => x"00000000",
 10258 => x"0000a2ac",
 10259 => x"0000a308",
 10260 => x"0000a364",
 10261 => x"00000000",
 10262 => x"00000000",
 10263 => x"00000000",
 10264 => x"00000000",
 10265 => x"00000000",
 10266 => x"00000000",
 10267 => x"00000000",
 10268 => x"00000000",
 10269 => x"00000000",
 10270 => x"00009e9c",
 10271 => x"00000000",
 10272 => x"00000000",
 10273 => x"00000000",
 10274 => x"00000000",
 10275 => x"00000000",
 10276 => x"00000000",
 10277 => x"00000000",
 10278 => x"00000000",
 10279 => x"00000000",
 10280 => x"00000000",
 10281 => x"00000000",
 10282 => x"00000000",
 10283 => x"00000000",
 10284 => x"00000000",
 10285 => x"00000000",
 10286 => x"00000000",
 10287 => x"00000000",
 10288 => x"00000000",
 10289 => x"00000000",
 10290 => x"00000000",
 10291 => x"00000000",
 10292 => x"00000000",
 10293 => x"00000000",
 10294 => x"00000000",
 10295 => x"00000000",
 10296 => x"00000000",
 10297 => x"00000000",
 10298 => x"00000000",
 10299 => x"00000001",
 10300 => x"330eabcd",
 10301 => x"1234e66d",
 10302 => x"deec0005",
 10303 => x"000b0000",
 10304 => x"00000000",
 10305 => x"00000000",
 10306 => x"00000000",
 10307 => x"00000000",
 10308 => x"00000000",
 10309 => x"00000000",
 10310 => x"00000000",
 10311 => x"00000000",
 10312 => x"00000000",
 10313 => x"00000000",
 10314 => x"00000000",
 10315 => x"00000000",
 10316 => x"00000000",
 10317 => x"00000000",
 10318 => x"00000000",
 10319 => x"00000000",
 10320 => x"00000000",
 10321 => x"00000000",
 10322 => x"00000000",
 10323 => x"00000000",
 10324 => x"00000000",
 10325 => x"00000000",
 10326 => x"00000000",
 10327 => x"00000000",
 10328 => x"00000000",
 10329 => x"00000000",
 10330 => x"00000000",
 10331 => x"00000000",
 10332 => x"00000000",
 10333 => x"00000000",
 10334 => x"00000000",
 10335 => x"00000000",
 10336 => x"00000000",
 10337 => x"00000000",
 10338 => x"00000000",
 10339 => x"00000000",
 10340 => x"00000000",
 10341 => x"00000000",
 10342 => x"00000000",
 10343 => x"00000000",
 10344 => x"00000000",
 10345 => x"00000000",
 10346 => x"00000000",
 10347 => x"00000000",
 10348 => x"00000000",
 10349 => x"00000000",
 10350 => x"00000000",
 10351 => x"00000000",
 10352 => x"00000000",
 10353 => x"00000000",
 10354 => x"00000000",
 10355 => x"00000000",
 10356 => x"00000000",
 10357 => x"00000000",
 10358 => x"00000000",
 10359 => x"00000000",
 10360 => x"00000000",
 10361 => x"00000000",
 10362 => x"00000000",
 10363 => x"00000000",
 10364 => x"00000000",
 10365 => x"00000000",
 10366 => x"00000000",
 10367 => x"00000000",
 10368 => x"00000000",
 10369 => x"00000000",
 10370 => x"00000000",
 10371 => x"00000000",
 10372 => x"00000000",
 10373 => x"00000000",
 10374 => x"00000000",
 10375 => x"00000000",
 10376 => x"00000000",
 10377 => x"00000000",
 10378 => x"00000000",
 10379 => x"00000000",
 10380 => x"00000000",
 10381 => x"00000000",
 10382 => x"00000000",
 10383 => x"00000000",
 10384 => x"00000000",
 10385 => x"00000000",
 10386 => x"00000000",
 10387 => x"00000000",
 10388 => x"00000000",
 10389 => x"00000000",
 10390 => x"00000000",
 10391 => x"00000000",
 10392 => x"00000000",
 10393 => x"00000000",
 10394 => x"00000000",
 10395 => x"00000000",
 10396 => x"00000000",
 10397 => x"00000000",
 10398 => x"00000000",
 10399 => x"00000000",
 10400 => x"00000000",
 10401 => x"00000000",
 10402 => x"00000000",
 10403 => x"00000000",
 10404 => x"00000000",
 10405 => x"00000000",
 10406 => x"00000000",
 10407 => x"00000000",
 10408 => x"00000000",
 10409 => x"00000000",
 10410 => x"00000000",
 10411 => x"00000000",
 10412 => x"00000000",
 10413 => x"00000000",
 10414 => x"00000000",
 10415 => x"00000000",
 10416 => x"00000000",
 10417 => x"00000000",
 10418 => x"00000000",
 10419 => x"00000000",
 10420 => x"00000000",
 10421 => x"00000000",
 10422 => x"00000000",
 10423 => x"00000000",
 10424 => x"00000000",
 10425 => x"00000000",
 10426 => x"00000000",
 10427 => x"00000000",
 10428 => x"00000000",
 10429 => x"00000000",
 10430 => x"00000000",
 10431 => x"00000000",
 10432 => x"00000000",
 10433 => x"00000000",
 10434 => x"00000000",
 10435 => x"00000000",
 10436 => x"00000000",
 10437 => x"00000000",
 10438 => x"00000000",
 10439 => x"00000000",
 10440 => x"00000000",
 10441 => x"00000000",
 10442 => x"00000000",
 10443 => x"00000000",
 10444 => x"00000000",
 10445 => x"00000000",
 10446 => x"00000000",
 10447 => x"00000000",
 10448 => x"00000000",
 10449 => x"00000000",
 10450 => x"00000000",
 10451 => x"00000000",
 10452 => x"00000000",
 10453 => x"00000000",
 10454 => x"00000000",
 10455 => x"00000000",
 10456 => x"00000000",
 10457 => x"00000000",
 10458 => x"00000000",
 10459 => x"00000000",
 10460 => x"00000000",
 10461 => x"00000000",
 10462 => x"00000000",
 10463 => x"00000000",
 10464 => x"00000000",
 10465 => x"00000000",
 10466 => x"00000000",
 10467 => x"00000000",
 10468 => x"00000000",
 10469 => x"00000000",
 10470 => x"00000000",
 10471 => x"00000000",
 10472 => x"00000000",
 10473 => x"00000000",
 10474 => x"00000000",
 10475 => x"00000000",
 10476 => x"00000000",
 10477 => x"00000000",
 10478 => x"00000000",
 10479 => x"00000000",
 10480 => x"43000000",
 10481 => x"00000000",
 10482 => x"00000000",
 10483 => x"00000000",
 10484 => x"00000000",
 10485 => x"00000000",
 10486 => x"00000001",
 10487 => x"00009ea0",
 10488 => x"00000000",
 10489 => x"00000000",
 10490 => x"00000000",
 10491 => x"00000000",
 10492 => x"00000000",
 10493 => x"00000000",
 10494 => x"00000000",
 10495 => x"00000000",
 10496 => x"00000000",
 10497 => x"00000000",
 10498 => x"00000000",
 10499 => x"00000000",
 10500 => x"ffffffff",
 10501 => x"00000000",
 10502 => x"00020000",
 10503 => x"00000000",
 10504 => x"00000000",
 10505 => x"0000a41c",
 10506 => x"0000a41c",
 10507 => x"0000a424",
 10508 => x"0000a424",
 10509 => x"0000a42c",
 10510 => x"0000a42c",
 10511 => x"0000a434",
 10512 => x"0000a434",
 10513 => x"0000a43c",
 10514 => x"0000a43c",
 10515 => x"0000a444",
 10516 => x"0000a444",
 10517 => x"0000a44c",
 10518 => x"0000a44c",
 10519 => x"0000a454",
 10520 => x"0000a454",
 10521 => x"0000a45c",
 10522 => x"0000a45c",
 10523 => x"0000a464",
 10524 => x"0000a464",
 10525 => x"0000a46c",
 10526 => x"0000a46c",
 10527 => x"0000a474",
 10528 => x"0000a474",
 10529 => x"0000a47c",
 10530 => x"0000a47c",
 10531 => x"0000a484",
 10532 => x"0000a484",
 10533 => x"0000a48c",
 10534 => x"0000a48c",
 10535 => x"0000a494",
 10536 => x"0000a494",
 10537 => x"0000a49c",
 10538 => x"0000a49c",
 10539 => x"0000a4a4",
 10540 => x"0000a4a4",
 10541 => x"0000a4ac",
 10542 => x"0000a4ac",
 10543 => x"0000a4b4",
 10544 => x"0000a4b4",
 10545 => x"0000a4bc",
 10546 => x"0000a4bc",
 10547 => x"0000a4c4",
 10548 => x"0000a4c4",
 10549 => x"0000a4cc",
 10550 => x"0000a4cc",
 10551 => x"0000a4d4",
 10552 => x"0000a4d4",
 10553 => x"0000a4dc",
 10554 => x"0000a4dc",
 10555 => x"0000a4e4",
 10556 => x"0000a4e4",
 10557 => x"0000a4ec",
 10558 => x"0000a4ec",
 10559 => x"0000a4f4",
 10560 => x"0000a4f4",
 10561 => x"0000a4fc",
 10562 => x"0000a4fc",
 10563 => x"0000a504",
 10564 => x"0000a504",
 10565 => x"0000a50c",
 10566 => x"0000a50c",
 10567 => x"0000a514",
 10568 => x"0000a514",
 10569 => x"0000a51c",
 10570 => x"0000a51c",
 10571 => x"0000a524",
 10572 => x"0000a524",
 10573 => x"0000a52c",
 10574 => x"0000a52c",
 10575 => x"0000a534",
 10576 => x"0000a534",
 10577 => x"0000a53c",
 10578 => x"0000a53c",
 10579 => x"0000a544",
 10580 => x"0000a544",
 10581 => x"0000a54c",
 10582 => x"0000a54c",
 10583 => x"0000a554",
 10584 => x"0000a554",
 10585 => x"0000a55c",
 10586 => x"0000a55c",
 10587 => x"0000a564",
 10588 => x"0000a564",
 10589 => x"0000a56c",
 10590 => x"0000a56c",
 10591 => x"0000a574",
 10592 => x"0000a574",
 10593 => x"0000a57c",
 10594 => x"0000a57c",
 10595 => x"0000a584",
 10596 => x"0000a584",
 10597 => x"0000a58c",
 10598 => x"0000a58c",
 10599 => x"0000a594",
 10600 => x"0000a594",
 10601 => x"0000a59c",
 10602 => x"0000a59c",
 10603 => x"0000a5a4",
 10604 => x"0000a5a4",
 10605 => x"0000a5ac",
 10606 => x"0000a5ac",
 10607 => x"0000a5b4",
 10608 => x"0000a5b4",
 10609 => x"0000a5bc",
 10610 => x"0000a5bc",
 10611 => x"0000a5c4",
 10612 => x"0000a5c4",
 10613 => x"0000a5cc",
 10614 => x"0000a5cc",
 10615 => x"0000a5d4",
 10616 => x"0000a5d4",
 10617 => x"0000a5dc",
 10618 => x"0000a5dc",
 10619 => x"0000a5e4",
 10620 => x"0000a5e4",
 10621 => x"0000a5ec",
 10622 => x"0000a5ec",
 10623 => x"0000a5f4",
 10624 => x"0000a5f4",
 10625 => x"0000a5fc",
 10626 => x"0000a5fc",
 10627 => x"0000a604",
 10628 => x"0000a604",
 10629 => x"0000a60c",
 10630 => x"0000a60c",
 10631 => x"0000a614",
 10632 => x"0000a614",
 10633 => x"0000a61c",
 10634 => x"0000a61c",
 10635 => x"0000a624",
 10636 => x"0000a624",
 10637 => x"0000a62c",
 10638 => x"0000a62c",
 10639 => x"0000a634",
 10640 => x"0000a634",
 10641 => x"0000a63c",
 10642 => x"0000a63c",
 10643 => x"0000a644",
 10644 => x"0000a644",
 10645 => x"0000a64c",
 10646 => x"0000a64c",
 10647 => x"0000a654",
 10648 => x"0000a654",
 10649 => x"0000a65c",
 10650 => x"0000a65c",
 10651 => x"0000a664",
 10652 => x"0000a664",
 10653 => x"0000a66c",
 10654 => x"0000a66c",
 10655 => x"0000a674",
 10656 => x"0000a674",
 10657 => x"0000a67c",
 10658 => x"0000a67c",
 10659 => x"0000a684",
 10660 => x"0000a684",
 10661 => x"0000a68c",
 10662 => x"0000a68c",
 10663 => x"0000a694",
 10664 => x"0000a694",
 10665 => x"0000a69c",
 10666 => x"0000a69c",
 10667 => x"0000a6a4",
 10668 => x"0000a6a4",
 10669 => x"0000a6ac",
 10670 => x"0000a6ac",
 10671 => x"0000a6b4",
 10672 => x"0000a6b4",
 10673 => x"0000a6bc",
 10674 => x"0000a6bc",
 10675 => x"0000a6c4",
 10676 => x"0000a6c4",
 10677 => x"0000a6cc",
 10678 => x"0000a6cc",
 10679 => x"0000a6d4",
 10680 => x"0000a6d4",
 10681 => x"0000a6dc",
 10682 => x"0000a6dc",
 10683 => x"0000a6e4",
 10684 => x"0000a6e4",
 10685 => x"0000a6ec",
 10686 => x"0000a6ec",
 10687 => x"0000a6f4",
 10688 => x"0000a6f4",
 10689 => x"0000a6fc",
 10690 => x"0000a6fc",
 10691 => x"0000a704",
 10692 => x"0000a704",
 10693 => x"0000a70c",
 10694 => x"0000a70c",
 10695 => x"0000a714",
 10696 => x"0000a714",
 10697 => x"0000a71c",
 10698 => x"0000a71c",
 10699 => x"0000a724",
 10700 => x"0000a724",
 10701 => x"0000a72c",
 10702 => x"0000a72c",
 10703 => x"0000a734",
 10704 => x"0000a734",
 10705 => x"0000a73c",
 10706 => x"0000a73c",
 10707 => x"0000a744",
 10708 => x"0000a744",
 10709 => x"0000a74c",
 10710 => x"0000a74c",
 10711 => x"0000a754",
 10712 => x"0000a754",
 10713 => x"0000a75c",
 10714 => x"0000a75c",
 10715 => x"0000a764",
 10716 => x"0000a764",
 10717 => x"0000a76c",
 10718 => x"0000a76c",
 10719 => x"0000a774",
 10720 => x"0000a774",
 10721 => x"0000a77c",
 10722 => x"0000a77c",
 10723 => x"0000a784",
 10724 => x"0000a784",
 10725 => x"0000a78c",
 10726 => x"0000a78c",
 10727 => x"0000a794",
 10728 => x"0000a794",
 10729 => x"0000a79c",
 10730 => x"0000a79c",
 10731 => x"0000a7a4",
 10732 => x"0000a7a4",
 10733 => x"0000a7ac",
 10734 => x"0000a7ac",
 10735 => x"0000a7b4",
 10736 => x"0000a7b4",
 10737 => x"0000a7bc",
 10738 => x"0000a7bc",
 10739 => x"0000a7c4",
 10740 => x"0000a7c4",
 10741 => x"0000a7cc",
 10742 => x"0000a7cc",
 10743 => x"0000a7d4",
 10744 => x"0000a7d4",
 10745 => x"0000a7dc",
 10746 => x"0000a7dc",
 10747 => x"0000a7e4",
 10748 => x"0000a7e4",
 10749 => x"0000a7ec",
 10750 => x"0000a7ec",
 10751 => x"0000a7f4",
 10752 => x"0000a7f4",
 10753 => x"0000a7fc",
 10754 => x"0000a7fc",
 10755 => x"0000a804",
 10756 => x"0000a804",
 10757 => x"0000a80c",
 10758 => x"0000a80c",
 10759 => x"0000a814",
 10760 => x"0000a814",
 10761 => x"0000a000",
 10762 => x"ffffffff",
 10763 => x"00000000",
 10764 => x"ffffffff",
 10765 => x"00000000",
 10766 => x"00000000",
  others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture rtl; -- Entity: SinglePortRAM

