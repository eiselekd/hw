../../nand/nand_parameters.vh