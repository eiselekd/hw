aldec/sim0/nand/nand_parameters.vh